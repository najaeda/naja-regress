module jpeg_rzs_clone_94(input clk, input ena, input rst, input deni, input dci,
 input [3:0] rleni, input [3:0] sizei, input [11:0] ampi, output deno, output dco, output [3:0] rleno,
 output [3:0] sizeo, output [11:0] ampo);
wire _000_;
wire _001_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _118_;
wire _119_;
wire \amp[0] ;
wire \amp[10] ;
wire \amp[11] ;
wire \amp[1] ;
wire \amp[2] ;
wire \amp[3] ;
wire \amp[4] ;
wire \amp[5] ;
wire \amp[6] ;
wire \amp[7] ;
wire \amp[8] ;
wire \amp[9] ;
wire den;
wire \rlen[0] ;
wire \rlen[1] ;
wire \rlen[2] ;
wire \rlen[3] ;
wire \size[0] ;
wire \size[1] ;
wire \size[2] ;
wire \size[3] ;
wire state;

NAND2_X1 _120_ (
  .A1(rleni[1]),
  .A2(rleni[0]),
  .ZN(_045_)
);

NAND2_X1 _121_ (
  .A1(rleni[3]),
  .A2(rleni[2]),
  .ZN(_046_)
);

NOR2_X1 _122_ (
  .A1(_045_),
  .A2(_046_),
  .ZN(_047_)
);

NOR2_X1 _123_ (
  .A1(sizei[1]),
  .A2(sizei[0]),
  .ZN(_048_)
);

NOR2_X1 _124_ (
  .A1(sizei[3]),
  .A2(sizei[2]),
  .ZN(_049_)
);

NAND3_X1 _125_ (
  .A1(_047_),
  .A2(_048_),
  .A3(_049_),
  .ZN(_050_)
);

BUF_X4 _126_ (
  .A(ena),
  .Z(_051_)
);

NAND2_X4 _127_ (
  .A1(deni),
  .A2(_051_),
  .ZN(_052_)
);

BUF_X8 _128_ (
  .A(_052_),
  .Z(_053_)
);

INV_X1 _129_ (
  .A(_053_),
  .ZN(_054_)
);

NAND2_X1 _130_ (
  .A1(_050_),
  .A2(_054_),
  .ZN(_055_)
);

INV_X1 _131_ (
  .A(state),
  .ZN(_056_)
);

NAND2_X1 _132_ (
  .A1(_056_),
  .A2(_051_),
  .ZN(_057_)
);

NAND3_X1 _133_ (
  .A1(_057_),
  .A2(_053_),
  .A3(den),
  .ZN(_058_)
);

NAND2_X1 _134_ (
  .A1(_055_),
  .A2(_058_),
  .ZN(_000_)
);

NOR2_X1 _135_ (
  .A1(_052_),
  .A2(_056_),
  .ZN(_059_)
);

NOR2_X1 _136_ (
  .A1(rleni[1]),
  .A2(rleni[0]),
  .ZN(_060_)
);

NOR2_X1 _137_ (
  .A1(rleni[3]),
  .A2(rleni[2]),
  .ZN(_061_)
);

INV_X1 _138_ (
  .A(dci),
  .ZN(_062_)
);

NAND3_X1 _139_ (
  .A1(_060_),
  .A2(_061_),
  .A3(_062_),
  .ZN(_063_)
);

NAND2_X1 _140_ (
  .A1(_048_),
  .A2(_049_),
  .ZN(_064_)
);

OAI21_X1 _141_ (
  .A(_059_),
  .B1(_063_),
  .B2(_064_),
  .ZN(_065_)
);

INV_X1 _142_ (
  .A(den),
  .ZN(_066_)
);

INV_X1 _143_ (
  .A(deno),
  .ZN(_067_)
);

OAI22_X1 _144_ (
  .A1(_057_),
  .A2(_066_),
  .B1(_067_),
  .B2(_051_),
  .ZN(_068_)
);

INV_X1 _145_ (
  .A(_068_),
  .ZN(_069_)
);

NAND2_X1 _146_ (
  .A1(_065_),
  .A2(_069_),
  .ZN(_001_)
);

BUF_X4 _147_ (
  .A(_051_),
  .Z(_070_)
);

BUF_X4 _150_ (
  .A(_051_),
  .Z(_072_)
);

MUX2_X1 _151_ (
  .A(rleno[0]),
  .B(\rlen[0] ),
  .S(_072_),
  .Z(_003_)
);

MUX2_X1 _152_ (
  .A(rleno[1]),
  .B(\rlen[1] ),
  .S(_070_),
  .Z(_004_)
);

MUX2_X1 _153_ (
  .A(rleno[2]),
  .B(\rlen[2] ),
  .S(_072_),
  .Z(_005_)
);

MUX2_X1 _154_ (
  .A(rleno[3]),
  .B(\rlen[3] ),
  .S(_070_),
  .Z(_006_)
);

MUX2_X1 _155_ (
  .A(sizeo[0]),
  .B(\size[0] ),
  .S(_072_),
  .Z(_007_)
);

MUX2_X1 _156_ (
  .A(sizeo[1]),
  .B(\size[1] ),
  .S(_051_),
  .Z(_008_)
);

MUX2_X1 _157_ (
  .A(sizeo[2]),
  .B(\size[2] ),
  .S(_051_),
  .Z(_009_)
);

MUX2_X1 _158_ (
  .A(sizeo[3]),
  .B(\size[3] ),
  .S(_070_),
  .Z(_010_)
);

MUX2_X1 _159_ (
  .A(ampo[0]),
  .B(\amp[0] ),
  .S(_072_),
  .Z(_011_)
);

MUX2_X1 _160_ (
  .A(ampo[1]),
  .B(\amp[1] ),
  .S(_072_),
  .Z(_012_)
);

MUX2_X1 _161_ (
  .A(ampo[2]),
  .B(\amp[2] ),
  .S(_070_),
  .Z(_013_)
);

MUX2_X1 _162_ (
  .A(ampo[3]),
  .B(\amp[3] ),
  .S(_072_),
  .Z(_014_)
);

MUX2_X1 _163_ (
  .A(ampo[4]),
  .B(\amp[4] ),
  .S(_070_),
  .Z(_015_)
);

MUX2_X1 _164_ (
  .A(ampo[5]),
  .B(\amp[5] ),
  .S(_072_),
  .Z(_016_)
);

MUX2_X1 _165_ (
  .A(ampo[6]),
  .B(\amp[6] ),
  .S(_070_),
  .Z(_017_)
);

MUX2_X1 _166_ (
  .A(ampo[7]),
  .B(\amp[7] ),
  .S(_072_),
  .Z(_018_)
);

MUX2_X1 _167_ (
  .A(ampo[8]),
  .B(\amp[8] ),
  .S(_072_),
  .Z(_019_)
);

MUX2_X1 _168_ (
  .A(ampo[9]),
  .B(\amp[9] ),
  .S(_070_),
  .Z(_020_)
);

MUX2_X1 _169_ (
  .A(ampo[10]),
  .B(\amp[10] ),
  .S(_072_),
  .Z(_021_)
);

MUX2_X1 _170_ (
  .A(ampo[11]),
  .B(\amp[11] ),
  .S(_070_),
  .Z(_022_)
);

MUX2_X1 _172_ (
  .A(sizei[0]),
  .B(\size[0] ),
  .S(_053_),
  .Z(_024_)
);

BUF_X8 _173_ (
  .A(_052_),
  .Z(_073_)
);

MUX2_X1 _174_ (
  .A(sizei[1]),
  .B(\size[1] ),
  .S(_073_),
  .Z(_025_)
);

MUX2_X1 _175_ (
  .A(sizei[2]),
  .B(\size[2] ),
  .S(_053_),
  .Z(_026_)
);

MUX2_X1 _176_ (
  .A(sizei[3]),
  .B(\size[3] ),
  .S(_053_),
  .Z(_027_)
);

MUX2_X1 _177_ (
  .A(rleni[0]),
  .B(\rlen[0] ),
  .S(_053_),
  .Z(_028_)
);

MUX2_X1 _178_ (
  .A(rleni[1]),
  .B(\rlen[1] ),
  .S(_053_),
  .Z(_029_)
);

MUX2_X1 _179_ (
  .A(rleni[2]),
  .B(\rlen[2] ),
  .S(_053_),
  .Z(_030_)
);

MUX2_X1 _180_ (
  .A(rleni[3]),
  .B(\rlen[3] ),
  .S(_073_),
  .Z(_031_)
);

MUX2_X1 _181_ (
  .A(ampi[0]),
  .B(\amp[0] ),
  .S(_073_),
  .Z(_032_)
);

MUX2_X1 _182_ (
  .A(ampi[1]),
  .B(\amp[1] ),
  .S(_073_),
  .Z(_033_)
);

MUX2_X1 _183_ (
  .A(ampi[2]),
  .B(\amp[2] ),
  .S(_073_),
  .Z(_034_)
);

MUX2_X1 _184_ (
  .A(ampi[3]),
  .B(\amp[3] ),
  .S(_052_),
  .Z(_035_)
);

MUX2_X1 _185_ (
  .A(ampi[4]),
  .B(\amp[4] ),
  .S(_073_),
  .Z(_036_)
);

MUX2_X1 _186_ (
  .A(ampi[5]),
  .B(\amp[5] ),
  .S(_073_),
  .Z(_037_)
);

MUX2_X1 _187_ (
  .A(ampi[6]),
  .B(\amp[6] ),
  .S(_073_),
  .Z(_038_)
);

MUX2_X1 _188_ (
  .A(ampi[7]),
  .B(\amp[7] ),
  .S(_073_),
  .Z(_039_)
);

MUX2_X1 _189_ (
  .A(ampi[8]),
  .B(\amp[8] ),
  .S(_073_),
  .Z(_040_)
);

MUX2_X1 _190_ (
  .A(ampi[9]),
  .B(\amp[9] ),
  .S(_052_),
  .Z(_041_)
);

MUX2_X1 _191_ (
  .A(ampi[10]),
  .B(\amp[10] ),
  .S(_052_),
  .Z(_042_)
);

MUX2_X1 _192_ (
  .A(ampi[11]),
  .B(\amp[11] ),
  .S(_052_),
  .Z(_043_)
);

NAND2_X1 _193_ (
  .A1(_053_),
  .A2(state),
  .ZN(_074_)
);

OAI21_X1 _194_ (
  .A(_074_),
  .B1(_050_),
  .B2(_053_),
  .ZN(_044_)
);

DFF_X1 \amp[0]$_DFFE_PP_  (
  .D(_032_),
  .CK(clk),
  .Q(\amp[0] ),
  .QN(_087_)
);

DFF_X1 \amp[10]$_DFFE_PP_  (
  .D(_042_),
  .CK(clk),
  .Q(\amp[10] ),
  .QN(_077_)
);

DFF_X1 \amp[11]$_DFFE_PP_  (
  .D(_043_),
  .CK(clk),
  .Q(\amp[11] ),
  .QN(_076_)
);

DFF_X1 \amp[1]$_DFFE_PP_  (
  .D(_033_),
  .CK(clk),
  .Q(\amp[1] ),
  .QN(_086_)
);

DFF_X1 \amp[2]$_DFFE_PP_  (
  .D(_034_),
  .CK(clk),
  .Q(\amp[2] ),
  .QN(_085_)
);

DFF_X1 \amp[3]$_DFFE_PP_  (
  .D(_035_),
  .CK(clk),
  .Q(\amp[3] ),
  .QN(_084_)
);

DFF_X1 \amp[4]$_DFFE_PP_  (
  .D(_036_),
  .CK(clk),
  .Q(\amp[4] ),
  .QN(_083_)
);

DFF_X1 \amp[5]$_DFFE_PP_  (
  .D(_037_),
  .CK(clk),
  .Q(\amp[5] ),
  .QN(_082_)
);

DFF_X1 \amp[6]$_DFFE_PP_  (
  .D(_038_),
  .CK(clk),
  .Q(\amp[6] ),
  .QN(_081_)
);

DFF_X1 \amp[7]$_DFFE_PP_  (
  .D(_039_),
  .CK(clk),
  .Q(\amp[7] ),
  .QN(_080_)
);

DFF_X1 \amp[8]$_DFFE_PP_  (
  .D(_040_),
  .CK(clk),
  .Q(\amp[8] ),
  .QN(_079_)
);

DFF_X1 \amp[9]$_DFFE_PP_  (
  .D(_041_),
  .CK(clk),
  .Q(\amp[9] ),
  .QN(_078_)
);

DFF_X1 \ampo[0]$_DFFE_PP_  (
  .D(_011_),
  .CK(clk),
  .Q(ampo[0]),
  .QN(_108_)
);

DFF_X1 \ampo[10]$_DFFE_PP_  (
  .D(_021_),
  .CK(clk),
  .Q(ampo[10]),
  .QN(_098_)
);

DFF_X1 \ampo[11]$_DFFE_PP_  (
  .D(_022_),
  .CK(clk),
  .Q(ampo[11]),
  .QN(_097_)
);

DFF_X1 \ampo[1]$_DFFE_PP_  (
  .D(_012_),
  .CK(clk),
  .Q(ampo[1]),
  .QN(_107_)
);

DFF_X1 \ampo[2]$_DFFE_PP_  (
  .D(_013_),
  .CK(clk),
  .Q(ampo[2]),
  .QN(_106_)
);

DFF_X1 \ampo[3]$_DFFE_PP_  (
  .D(_014_),
  .CK(clk),
  .Q(ampo[3]),
  .QN(_105_)
);

DFF_X1 \ampo[4]$_DFFE_PP_  (
  .D(_015_),
  .CK(clk),
  .Q(ampo[4]),
  .QN(_104_)
);

DFF_X1 \ampo[5]$_DFFE_PP_  (
  .D(_016_),
  .CK(clk),
  .Q(ampo[5]),
  .QN(_103_)
);

DFF_X1 \ampo[6]$_DFFE_PP_  (
  .D(_017_),
  .CK(clk),
  .Q(ampo[6]),
  .QN(_102_)
);

DFF_X1 \ampo[7]$_DFFE_PP_  (
  .D(_018_),
  .CK(clk),
  .Q(ampo[7]),
  .QN(_101_)
);

DFF_X1 \ampo[8]$_DFFE_PP_  (
  .D(_019_),
  .CK(clk),
  .Q(ampo[8]),
  .QN(_100_)
);

DFF_X1 \ampo[9]$_DFFE_PP_  (
  .D(_020_),
  .CK(clk),
  .Q(ampo[9]),
  .QN(_099_)
);

DFFR_X1 den$_DFFE_PN0P_ (
  .D(_000_),
  .RN(rst),
  .CK(clk),
  .Q(den),
  .QN(_119_)
);

DFFR_X1 deno$_DFFE_PN0P_ (
  .D(_001_),
  .RN(rst),
  .CK(clk),
  .Q(deno),
  .QN(_118_)
);

DFF_X1 \rlen[0]$_DFFE_PP_  (
  .D(_028_),
  .CK(clk),
  .Q(\rlen[0] ),
  .QN(_091_)
);

DFF_X1 \rlen[1]$_DFFE_PP_  (
  .D(_029_),
  .CK(clk),
  .Q(\rlen[1] ),
  .QN(_090_)
);

DFF_X1 \rlen[2]$_DFFE_PP_  (
  .D(_030_),
  .CK(clk),
  .Q(\rlen[2] ),
  .QN(_089_)
);

DFF_X1 \rlen[3]$_DFFE_PP_  (
  .D(_031_),
  .CK(clk),
  .Q(\rlen[3] ),
  .QN(_088_)
);

DFF_X1 \rleno[0]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(rleno[0]),
  .QN(_116_)
);

DFF_X1 \rleno[1]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(rleno[1]),
  .QN(_115_)
);

DFF_X1 \rleno[2]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(rleno[2]),
  .QN(_114_)
);

DFF_X1 \rleno[3]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(rleno[3]),
  .QN(_113_)
);

DFF_X1 \size[0]$_DFFE_PP_  (
  .D(_024_),
  .CK(clk),
  .Q(\size[0] ),
  .QN(_095_)
);

DFF_X1 \size[1]$_DFFE_PP_  (
  .D(_025_),
  .CK(clk),
  .Q(\size[1] ),
  .QN(_094_)
);

DFF_X1 \size[2]$_DFFE_PP_  (
  .D(_026_),
  .CK(clk),
  .Q(\size[2] ),
  .QN(_093_)
);

DFF_X1 \size[3]$_DFFE_PP_  (
  .D(_027_),
  .CK(clk),
  .Q(\size[3] ),
  .QN(_092_)
);

DFF_X1 \sizeo[0]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(sizeo[0]),
  .QN(_112_)
);

DFF_X1 \sizeo[1]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(sizeo[1]),
  .QN(_111_)
);

DFF_X1 \sizeo[2]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(sizeo[2]),
  .QN(_110_)
);

DFF_X1 \sizeo[3]$_DFFE_PP_  (
  .D(_010_),
  .CK(clk),
  .Q(sizeo[3]),
  .QN(_109_)
);

DFFR_X1 state$_DFFE_PN0P_ (
  .D(_044_),
  .RN(rst),
  .CK(clk),
  .Q(state),
  .QN(_075_)
);
endmodule //jpeg_rzs_clone_94

module \$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 (input clk,
 input ena, input dclr, input [7:0] din, input [10:0] coef, output [21:0] result);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire _0032_;
wire _0033_;
wire _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire _0066_;
wire _0067_;
wire _0068_;
wire _0069_;
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0333_;
wire _0339_;
wire _0341_;
wire _0348_;
wire _0354_;
wire _0355_;
wire _0367_;
wire _0368_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
wire _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
wire _0444_;
wire _0445_;
wire _0446_;
wire _0447_;
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0518_;
wire _0519_;
wire _0521_;
wire _0522_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire _0658_;
wire _0659_;
wire _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire _0673_;
wire _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire _0679_;
wire _0680_;
wire _0684_;
wire _0685_;
wire _0689_;
wire _0690_;
wire _0692_;
wire _0693_;
wire _0697_;
wire _0698_;
wire _0699_;
wire _0700_;
wire _0701_;
wire _0702_;
wire _0706_;
wire _0707_;
wire _0711_;
wire _0712_;
wire _0713_;
wire _0714_;
wire _0715_;
wire _0716_;
wire _0717_;
wire _0718_;
wire _0719_;
wire _0723_;
wire _0724_;
wire _0728_;
wire _0729_;
wire _0730_;
wire _0731_;
wire _0732_;
wire _0733_;
wire _0734_;
wire _0735_;
wire _0738_;
wire _0739_;
wire _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0751_;
wire _0752_;
wire _0756_;
wire _0757_;
wire _0761_;
wire _0762_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire _0780_;
wire _0781_;
wire _0782_;
wire _0783_;
wire _0784_;
wire _0785_;
wire _0786_;
wire _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire _0796_;
wire _0798_;
wire _0799_;
wire _0803_;
wire _0804_;
wire _0805_;
wire _0806_;
wire _0809_;
wire _0810_;
wire _0811_;
wire _0812_;
wire _0813_;
wire _0814_;
wire _0815_;
wire _0816_;
wire _0817_;
wire _0818_;
wire _0819_;
wire _0820_;
wire _0823_;
wire _0824_;
wire _0825_;
wire _0829_;
wire _0830_;
wire _0831_;
wire _0832_;
wire _0835_;
wire _0836_;
wire _0837_;
wire _0838_;
wire _0839_;
wire _0840_;
wire _0841_;
wire _0842_;
wire _0843_;
wire _0844_;
wire _0845_;
wire _0846_;
wire _0847_;
wire _0848_;
wire _0849_;
wire _0850_;
wire _0851_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0860_;
wire _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0867_;
wire _0868_;
wire _0869_;
wire _0870_;
wire _0871_;
wire _0872_;
wire _0874_;
wire _0875_;
wire _0876_;
wire _0877_;
wire _0878_;
wire _0879_;
wire _0880_;
wire _0881_;
wire _0883_;
wire _0884_;
wire _0886_;
wire _0888_;
wire _0889_;
wire _0890_;
wire _0891_;
wire _0892_;
wire _0893_;
wire _0896_;
wire _0897_;
wire _0898_;
wire _0899_;
wire _0900_;
wire _0901_;
wire _0902_;
wire _0903_;
wire _0904_;
wire _0905_;
wire _0906_;
wire _0907_;
wire _0908_;
wire _0909_;
wire _0910_;
wire _0911_;
wire _0912_;
wire _0913_;
wire _0914_;
wire _0915_;
wire _0916_;
wire _0917_;
wire _0918_;
wire _0921_;
wire _0922_;
wire _0923_;
wire _0924_;
wire _0925_;
wire _0926_;
wire _0929_;
wire _0930_;
wire _0931_;
wire _0932_;
wire _0933_;
wire _0934_;
wire _0935_;
wire _0936_;
wire _0937_;
wire _0938_;
wire _0939_;
wire _0940_;
wire _0941_;
wire _0942_;
wire _0943_;
wire _0944_;
wire _0945_;
wire _0946_;
wire _0947_;
wire _0948_;
wire _0949_;
wire _0950_;
wire _0954_;
wire _0955_;
wire _0956_;
wire _0957_;
wire _0958_;
wire _0959_;
wire _0961_;
wire _0962_;
wire _0963_;
wire _0964_;
wire _0965_;
wire _0966_;
wire _0967_;
wire _0968_;
wire _0969_;
wire _0970_;
wire _0971_;
wire _0972_;
wire _0973_;
wire _0974_;
wire _0975_;
wire _0976_;
wire _0977_;
wire _0978_;
wire _0979_;
wire _0980_;
wire _0981_;
wire _0982_;
wire _0983_;
wire _0984_;
wire _0985_;
wire _0987_;
wire _0988_;
wire _0989_;
wire _0990_;
wire _0991_;
wire _0993_;
wire _0994_;
wire _0995_;
wire _0996_;
wire _0997_;
wire _0998_;
wire _0999_;
wire _1000_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire \ext_mult_res[0] ;
wire \ext_mult_res[10] ;
wire \ext_mult_res[11] ;
wire \ext_mult_res[12] ;
wire \ext_mult_res[13] ;
wire \ext_mult_res[14] ;
wire \ext_mult_res[15] ;
wire \ext_mult_res[16] ;
wire \ext_mult_res[17] ;
wire \ext_mult_res[18] ;
wire \ext_mult_res[1] ;
wire \ext_mult_res[2] ;
wire \ext_mult_res[3] ;
wire \ext_mult_res[4] ;
wire \ext_mult_res[5] ;
wire \ext_mult_res[6] ;
wire \ext_mult_res[7] ;
wire \ext_mult_res[8] ;
wire \ext_mult_res[9] ;
wire \logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ;
wire \logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ;

BUF_X1 _1235_ (
  .A(din[0]),
  .Z(_0326_)
);

BUF_X1 _1245_ (
  .A(din[1]),
  .Z(_0333_)
);

BUF_X1 _1255_ (
  .A(din[2]),
  .Z(_0339_)
);

BUF_X1 _1258_ (
  .A(din[3]),
  .Z(_0341_)
);

BUF_X1 _1279_ (
  .A(din[6]),
  .Z(_0348_)
);

BUF_X1 _1292_ (
  .A(din[4]),
  .Z(_0354_)
);

BUF_X1 _1294_ (
  .A(din[5]),
  .Z(_0355_)
);

INV_X1 _1342_ (
  .A(_1177_),
  .ZN(_0792_)
);

INV_X1 _1360_ (
  .A(_0993_),
  .ZN(_1022_)
);

INV_X1 _1365_ (
  .A(_0987_),
  .ZN(_1027_)
);

INV_X1 _1366_ (
  .A(_0874_),
  .ZN(_0905_)
);

INV_X1 _1368_ (
  .A(_0785_),
  .ZN(_0786_)
);

INV_X1 _1370_ (
  .A(_0875_),
  .ZN(_0969_)
);

INV_X1 _1374_ (
  .A(_0903_),
  .ZN(_0904_)
);

INV_X1 _1376_ (
  .A(_0936_),
  .ZN(_0938_)
);

INV_X1 _1377_ (
  .A(_0968_),
  .ZN(_0970_)
);

INV_X1 _1378_ (
  .A(_1088_),
  .ZN(_0678_)
);

INV_X1 _1381_ (
  .A(_1152_),
  .ZN(_0787_)
);

INV_X1 _1382_ (
  .A(_1186_),
  .ZN(_0879_)
);

INV_X1 _1383_ (
  .A(_1193_),
  .ZN(_0916_)
);

INV_X1 _1385_ (
  .A(_1029_),
  .ZN(_1067_)
);

INV_X1 _1386_ (
  .A(_0752_),
  .ZN(_0775_)
);

INV_X1 _1387_ (
  .A(_0769_),
  .ZN(_0771_)
);

INV_X1 _1388_ (
  .A(_0856_),
  .ZN(_0862_)
);

INV_X1 _1389_ (
  .A(_0884_),
  .ZN(_0890_)
);

INV_X1 _1390_ (
  .A(_0912_),
  .ZN(_0913_)
);

INV_X1 _1391_ (
  .A(_0950_),
  .ZN(_1204_)
);

INV_X1 _1392_ (
  .A(_0955_),
  .ZN(_0956_)
);

INV_X1 _1393_ (
  .A(_0985_),
  .ZN(_1211_)
);

INV_X1 _1394_ (
  .A(_0988_),
  .ZN(_0989_)
);

INV_X1 _1395_ (
  .A(_1026_),
  .ZN(_1028_)
);

INV_X1 _1396_ (
  .A(_1037_),
  .ZN(_1038_)
);

INV_X1 _1397_ (
  .A(_1056_),
  .ZN(_1057_)
);

INV_X1 _1398_ (
  .A(_1079_),
  .ZN(_1080_)
);

INV_X1 _1399_ (
  .A(_0689_),
  .ZN(_0699_)
);

INV_X1 _1400_ (
  .A(_0751_),
  .ZN(_0745_)
);

INV_X1 _1401_ (
  .A(_0776_),
  .ZN(_0770_)
);

INV_X1 _1402_ (
  .A(_0855_),
  .ZN(_0891_)
);

INV_X1 _1403_ (
  .A(_0883_),
  .ZN(_0924_)
);

INV_X1 _1404_ (
  .A(_0954_),
  .ZN(_0996_)
);

INV_X1 _1405_ (
  .A(_1007_),
  .ZN(_1039_)
);

INV_X1 _1406_ (
  .A(_1025_),
  .ZN(_1058_)
);

INV_X1 _1407_ (
  .A(_0702_),
  .ZN(_1141_)
);

INV_X1 _1408_ (
  .A(_0714_),
  .ZN(_0715_)
);

INV_X1 _1409_ (
  .A(_0711_),
  .ZN(_1150_)
);

INV_X1 _1410_ (
  .A(_0734_),
  .ZN(_1154_)
);

INV_X1 _1413_ (
  .A(_0723_),
  .ZN(_0774_)
);

INV_X1 _1414_ (
  .A(_0756_),
  .ZN(_0765_)
);

INV_X1 _1415_ (
  .A(_0728_),
  .ZN(_1163_)
);

INV_X1 _1416_ (
  .A(_0773_),
  .ZN(_0778_)
);

INV_X1 _1417_ (
  .A(_0789_),
  .ZN(_1171_)
);

INV_X1 _1418_ (
  .A(_0743_),
  .ZN(_0811_)
);

INV_X1 _1419_ (
  .A(_0820_),
  .ZN(_1179_)
);

INV_X1 _1420_ (
  .A(_0836_),
  .ZN(_0838_)
);

INV_X1 _1421_ (
  .A(_0809_),
  .ZN(_0837_)
);

INV_X1 _1422_ (
  .A(_0846_),
  .ZN(_0848_)
);

INV_X1 _1423_ (
  .A(_0869_),
  .ZN(_0908_)
);

INV_X1 _1424_ (
  .A(_0880_),
  .ZN(_1199_)
);

INV_X1 _1425_ (
  .A(_0946_),
  .ZN(_0947_)
);

INV_X1 _1426_ (
  .A(_0931_),
  .ZN(_0974_)
);

INV_X1 _1427_ (
  .A(_0945_),
  .ZN(_0982_)
);

INV_X1 _1428_ (
  .A(_0943_),
  .ZN(_1210_)
);

INV_X1 _1429_ (
  .A(_0991_),
  .ZN(_1216_)
);

INV_X1 _1430_ (
  .A(_0963_),
  .ZN(_1009_)
);

INV_X1 _1431_ (
  .A(_1017_),
  .ZN(_1018_)
);

INV_X1 _1432_ (
  .A(_0990_),
  .ZN(_1222_)
);

INV_X1 _1433_ (
  .A(_1046_),
  .ZN(_1047_)
);

INV_X1 _1434_ (
  .A(_1040_),
  .ZN(_1075_)
);

INV_X1 _1435_ (
  .A(_1082_),
  .ZN(_1083_)
);

INV_X1 _1436_ (
  .A(_0701_),
  .ZN(_0716_)
);

INV_X1 _1437_ (
  .A(_0762_),
  .ZN(_0766_)
);

INV_X1 _1438_ (
  .A(_0783_),
  .ZN(_0779_)
);

INV_X1 _1439_ (
  .A(_0788_),
  .ZN(_1165_)
);

INV_X1 _1440_ (
  .A(_0810_),
  .ZN(_0812_)
);

INV_X1 _1441_ (
  .A(_0761_),
  .ZN(_0813_)
);

INV_X1 _1442_ (
  .A(_0803_),
  .ZN(_0839_)
);

INV_X1 _1443_ (
  .A(_0819_),
  .ZN(_0849_)
);

INV_X1 _1444_ (
  .A(_0907_),
  .ZN(_0909_)
);

INV_X1 _1445_ (
  .A(_0914_),
  .ZN(_0948_)
);

INV_X1 _1446_ (
  .A(_0917_),
  .ZN(_1205_)
);

INV_X1 _1447_ (
  .A(_0935_),
  .ZN(_0973_)
);

INV_X1 _1448_ (
  .A(_0972_),
  .ZN(_0975_)
);

INV_X1 _1449_ (
  .A(_0939_),
  .ZN(_0976_)
);

INV_X1 _1450_ (
  .A(_0980_),
  .ZN(_0983_)
);

INV_X1 _1451_ (
  .A(_0967_),
  .ZN(_1006_)
);

INV_X1 _1452_ (
  .A(_0971_),
  .ZN(_1010_)
);

INV_X1 _1453_ (
  .A(_0902_),
  .ZN(_0942_)
);

INV_X1 _1454_ (
  .A(_1016_),
  .ZN(_1048_)
);

INV_X1 _1455_ (
  .A(_1045_),
  .ZN(_1084_)
);

INV_X1 _1456_ (
  .A(_1153_),
  .ZN(_0732_)
);

INV_X1 _1457_ (
  .A(_1170_),
  .ZN(_0790_)
);

INV_X1 _1458_ (
  .A(_1178_),
  .ZN(_0818_)
);

INV_X1 _1459_ (
  .A(_1187_),
  .ZN(_0844_)
);

INV_X1 _1460_ (
  .A(_1194_),
  .ZN(_0876_)
);

INV_X1 _1461_ (
  .A(_1219_),
  .ZN(_1015_)
);

INV_X1 _1462_ (
  .A(_1228_),
  .ZN(_1044_)
);

INV_X1 _1463_ (
  .A(_1140_),
  .ZN(_0700_)
);

INV_X1 _1464_ (
  .A(_1164_),
  .ZN(_0784_)
);

INV_X1 _1465_ (
  .A(_0941_),
  .ZN(_0937_)
);

INV_X1 _1466_ (
  .A(_1173_),
  .ZN(_0791_)
);

BUF_X1 _1467_ (
  .A(ena),
  .Z(_0367_)
);

BUF_X1 _1468_ (
  .A(_0367_),
  .Z(_0368_)
);

INV_X1 _1470_ (
  .A(\ext_mult_res[0] ),
  .ZN(_0370_)
);

BUF_X1 _1471_ (
  .A(_0367_),
  .Z(_0371_)
);

BUF_X1 _1472_ (
  .A(_0371_),
  .Z(_0372_)
);

BUF_X1 _1474_ (
  .A(_0367_),
  .Z(_0373_)
);

MUX2_X1 _1475_ (
  .A(\ext_mult_res[1] ),
  .B(_1133_),
  .S(_0373_),
  .Z(_0001_)
);

BUF_X4 _1476_ (
  .A(_0371_),
  .Z(_0374_)
);

NAND2_X1 _1477_ (
  .A1(_0374_),
  .A2(_1135_),
  .ZN(_0375_)
);

INV_X1 _1478_ (
  .A(\ext_mult_res[2] ),
  .ZN(_0376_)
);

OAI21_X1 _1479_ (
  .A(_0375_),
  .B1(_0376_),
  .B2(_0372_),
  .ZN(_0002_)
);

NAND2_X1 _1480_ (
  .A1(_0374_),
  .A2(_1137_),
  .ZN(_0377_)
);

INV_X1 _1481_ (
  .A(\ext_mult_res[3] ),
  .ZN(_0378_)
);

OAI21_X1 _1482_ (
  .A(_0377_),
  .B1(_0378_),
  .B2(_0372_),
  .ZN(_0003_)
);

NAND2_X1 _1483_ (
  .A1(_0374_),
  .A2(_1145_),
  .ZN(_0379_)
);

INV_X1 _1484_ (
  .A(\ext_mult_res[4] ),
  .ZN(_0380_)
);

OAI21_X1 _1485_ (
  .A(_0379_),
  .B1(_0380_),
  .B2(_0372_),
  .ZN(_0004_)
);

MUX2_X1 _1486_ (
  .A(\ext_mult_res[5] ),
  .B(_1149_),
  .S(_0373_),
  .Z(_0005_)
);

NAND2_X1 _1487_ (
  .A1(_0372_),
  .A2(_1160_),
  .ZN(_0381_)
);

INV_X1 _1488_ (
  .A(\ext_mult_res[6] ),
  .ZN(_0382_)
);

OAI21_X1 _1489_ (
  .A(_0381_),
  .B1(_0382_),
  .B2(_0372_),
  .ZN(_0006_)
);

NAND2_X1 _1490_ (
  .A1(_0374_),
  .A2(_1234_),
  .ZN(_0383_)
);

INV_X1 _1491_ (
  .A(\ext_mult_res[7] ),
  .ZN(_0384_)
);

OAI21_X1 _1492_ (
  .A(_0383_),
  .B1(_0384_),
  .B2(_0372_),
  .ZN(_0007_)
);

INV_X1 _1493_ (
  .A(_0367_),
  .ZN(_0385_)
);

NAND2_X1 _1494_ (
  .A1(_0385_),
  .A2(\ext_mult_res[8] ),
  .ZN(_0386_)
);

BUF_X1 _1495_ (
  .A(_0385_),
  .Z(_0387_)
);

OAI21_X1 _1496_ (
  .A(_0386_),
  .B1(_0794_),
  .B2(_0387_),
  .ZN(_0008_)
);

INV_X1 _1497_ (
  .A(_0793_),
  .ZN(_0388_)
);

NAND2_X1 _1498_ (
  .A1(_0388_),
  .A2(_1185_),
  .ZN(_0389_)
);

INV_X1 _1499_ (
  .A(_1185_),
  .ZN(_0390_)
);

NAND2_X1 _1500_ (
  .A1(_0390_),
  .A2(_0793_),
  .ZN(_0391_)
);

NAND3_X1 _1501_ (
  .A1(_0389_),
  .A2(_0391_),
  .A3(_0374_),
  .ZN(_0392_)
);

INV_X1 _1502_ (
  .A(\ext_mult_res[9] ),
  .ZN(_0393_)
);

OAI21_X1 _1503_ (
  .A(_0392_),
  .B1(_0393_),
  .B2(_0372_),
  .ZN(_0009_)
);

NOR2_X1 _1504_ (
  .A1(\ext_mult_res[10] ),
  .A2(_0373_),
  .ZN(_0394_)
);

INV_X1 _1505_ (
  .A(_1184_),
  .ZN(_0395_)
);

INV_X1 _1506_ (
  .A(_1174_),
  .ZN(_0396_)
);

OAI21_X1 _1507_ (
  .A(_0395_),
  .B1(_0390_),
  .B2(_0396_),
  .ZN(_0397_)
);

INV_X1 _1508_ (
  .A(_0397_),
  .ZN(_0398_)
);

NAND2_X1 _1509_ (
  .A1(_1185_),
  .A2(_1175_),
  .ZN(_0399_)
);

OAI21_X1 _1510_ (
  .A(_0398_),
  .B1(_0792_),
  .B2(_0399_),
  .ZN(_0400_)
);

BUF_X1 _1511_ (
  .A(_1191_),
  .Z(_0401_)
);

XNOR2_X1 _1512_ (
  .A(_0400_),
  .B(_0401_),
  .ZN(_0402_)
);

BUF_X1 _1513_ (
  .A(_0371_),
  .Z(_0403_)
);

AOI21_X1 _1514_ (
  .A(_0394_),
  .B1(_0402_),
  .B2(_0403_),
  .ZN(_0010_)
);

NOR2_X1 _1515_ (
  .A1(\ext_mult_res[11] ),
  .A2(_0373_),
  .ZN(_0404_)
);

INV_X1 _1516_ (
  .A(_1190_),
  .ZN(_0405_)
);

INV_X1 _1517_ (
  .A(_0401_),
  .ZN(_0406_)
);

OAI21_X1 _1518_ (
  .A(_0405_),
  .B1(_0406_),
  .B2(_0395_),
  .ZN(_0407_)
);

NAND2_X1 _1519_ (
  .A1(_1185_),
  .A2(_0401_),
  .ZN(_0408_)
);

INV_X1 _1520_ (
  .A(_0408_),
  .ZN(_0409_)
);

AOI21_X1 _1521_ (
  .A(_0407_),
  .B1(_0409_),
  .B2(_0388_),
  .ZN(_0410_)
);

INV_X1 _1522_ (
  .A(_1198_),
  .ZN(_0411_)
);

XNOR2_X1 _1523_ (
  .A(_0410_),
  .B(_0411_),
  .ZN(_0412_)
);

AOI21_X1 _1524_ (
  .A(_0404_),
  .B1(_0412_),
  .B2(_0403_),
  .ZN(_0011_)
);

NOR2_X1 _1525_ (
  .A1(\ext_mult_res[12] ),
  .A2(_0373_),
  .ZN(_0413_)
);

INV_X1 _1526_ (
  .A(_1197_),
  .ZN(_0414_)
);

OAI21_X1 _1527_ (
  .A(_0414_),
  .B1(_0411_),
  .B2(_0405_),
  .ZN(_0415_)
);

INV_X1 _1528_ (
  .A(_0415_),
  .ZN(_0416_)
);

NAND2_X1 _1529_ (
  .A1(_0401_),
  .A2(_1198_),
  .ZN(_0417_)
);

OAI21_X1 _1530_ (
  .A(_0416_),
  .B1(_0398_),
  .B2(_0417_),
  .ZN(_0418_)
);

NOR2_X1 _1531_ (
  .A1(_0399_),
  .A2(_0417_),
  .ZN(_0419_)
);

AOI21_X1 _1532_ (
  .A(_0418_),
  .B1(_0419_),
  .B2(_1177_),
  .ZN(_0420_)
);

INV_X1 _1533_ (
  .A(_1203_),
  .ZN(_0421_)
);

XNOR2_X1 _1534_ (
  .A(_0420_),
  .B(_0421_),
  .ZN(_0422_)
);

AOI21_X1 _1535_ (
  .A(_0413_),
  .B1(_0422_),
  .B2(_0403_),
  .ZN(_0012_)
);

NOR2_X1 _1536_ (
  .A1(\ext_mult_res[13] ),
  .A2(_0373_),
  .ZN(_0423_)
);

INV_X1 _1537_ (
  .A(_1202_),
  .ZN(_0424_)
);

OAI21_X1 _1538_ (
  .A(_0424_),
  .B1(_0421_),
  .B2(_0414_),
  .ZN(_0425_)
);

INV_X1 _1539_ (
  .A(_0425_),
  .ZN(_0426_)
);

INV_X1 _1540_ (
  .A(_0407_),
  .ZN(_0427_)
);

NAND2_X1 _1541_ (
  .A1(_1198_),
  .A2(_1203_),
  .ZN(_0428_)
);

OAI21_X1 _1542_ (
  .A(_0426_),
  .B1(_0427_),
  .B2(_0428_),
  .ZN(_0429_)
);

NOR2_X1 _1543_ (
  .A1(_0408_),
  .A2(_0428_),
  .ZN(_0430_)
);

AOI21_X1 _1544_ (
  .A(_0429_),
  .B1(_0430_),
  .B2(_0388_),
  .ZN(_0431_)
);

INV_X1 _1545_ (
  .A(_1209_),
  .ZN(_0432_)
);

XNOR2_X1 _1546_ (
  .A(_0431_),
  .B(_0432_),
  .ZN(_0433_)
);

AOI21_X1 _1547_ (
  .A(_0423_),
  .B1(_0433_),
  .B2(_0403_),
  .ZN(_0013_)
);

NOR2_X1 _1548_ (
  .A1(\ext_mult_res[14] ),
  .A2(_0373_),
  .ZN(_0434_)
);

INV_X1 _1549_ (
  .A(_1208_),
  .ZN(_0435_)
);

OAI21_X1 _1550_ (
  .A(_0435_),
  .B1(_0432_),
  .B2(_0424_),
  .ZN(_0436_)
);

INV_X1 _1551_ (
  .A(_0436_),
  .ZN(_0437_)
);

NAND2_X1 _1552_ (
  .A1(_1203_),
  .A2(_1209_),
  .ZN(_0438_)
);

OAI21_X1 _1553_ (
  .A(_0437_),
  .B1(_0416_),
  .B2(_0438_),
  .ZN(_0439_)
);

NOR2_X1 _1554_ (
  .A1(_0417_),
  .A2(_0438_),
  .ZN(_0440_)
);

AOI21_X1 _1555_ (
  .A(_0439_),
  .B1(_0440_),
  .B2(_0400_),
  .ZN(_0441_)
);

INV_X1 _1556_ (
  .A(_1215_),
  .ZN(_0442_)
);

XNOR2_X1 _1557_ (
  .A(_0441_),
  .B(_0442_),
  .ZN(_0443_)
);

AOI21_X1 _1558_ (
  .A(_0434_),
  .B1(_0443_),
  .B2(_0403_),
  .ZN(_0014_)
);

NAND2_X1 _1559_ (
  .A1(_1209_),
  .A2(_1215_),
  .ZN(_0444_)
);

NOR3_X1 _1560_ (
  .A1(_0410_),
  .A2(_0428_),
  .A3(_0444_),
  .ZN(_0445_)
);

INV_X1 _1561_ (
  .A(_1214_),
  .ZN(_0446_)
);

OAI21_X1 _1562_ (
  .A(_0446_),
  .B1(_0442_),
  .B2(_0435_),
  .ZN(_0447_)
);

INV_X1 _1563_ (
  .A(_0447_),
  .ZN(_0448_)
);

OAI21_X1 _1564_ (
  .A(_0448_),
  .B1(_0426_),
  .B2(_0444_),
  .ZN(_0449_)
);

OR2_X1 _1565_ (
  .A1(_0445_),
  .A2(_0449_),
  .ZN(_0450_)
);

BUF_X1 _1566_ (
  .A(_1221_),
  .Z(_0451_)
);

OR2_X1 _1567_ (
  .A1(_0450_),
  .A2(_0451_),
  .ZN(_0452_)
);

NAND2_X1 _1568_ (
  .A1(_0450_),
  .A2(_0451_),
  .ZN(_0453_)
);

NAND3_X1 _1569_ (
  .A1(_0452_),
  .A2(_0374_),
  .A3(_0453_),
  .ZN(_0454_)
);

INV_X1 _1570_ (
  .A(\ext_mult_res[15] ),
  .ZN(_0455_)
);

OAI21_X1 _1571_ (
  .A(_0454_),
  .B1(_0455_),
  .B2(_0372_),
  .ZN(_0015_)
);

NOR2_X1 _1572_ (
  .A1(\ext_mult_res[16] ),
  .A2(_0373_),
  .ZN(_0456_)
);

INV_X1 _1573_ (
  .A(_1220_),
  .ZN(_0457_)
);

INV_X1 _1574_ (
  .A(_0451_),
  .ZN(_0458_)
);

OAI21_X1 _1575_ (
  .A(_0457_),
  .B1(_0458_),
  .B2(_0446_),
  .ZN(_0459_)
);

INV_X1 _1576_ (
  .A(_0459_),
  .ZN(_0460_)
);

NAND2_X1 _1577_ (
  .A1(_1215_),
  .A2(_0451_),
  .ZN(_0461_)
);

OAI21_X1 _1578_ (
  .A(_0460_),
  .B1(_0437_),
  .B2(_0461_),
  .ZN(_0462_)
);

NOR2_X1 _1579_ (
  .A1(_0438_),
  .A2(_0461_),
  .ZN(_0463_)
);

AOI21_X1 _1580_ (
  .A(_0462_),
  .B1(_0463_),
  .B2(_0418_),
  .ZN(_0464_)
);

NAND3_X1 _1581_ (
  .A1(_0419_),
  .A2(_0463_),
  .A3(_1177_),
  .ZN(_0465_)
);

NAND2_X1 _1582_ (
  .A1(_0464_),
  .A2(_0465_),
  .ZN(_0466_)
);

BUF_X1 _1583_ (
  .A(_1230_),
  .Z(_0467_)
);

XNOR2_X1 _1584_ (
  .A(_0466_),
  .B(_0467_),
  .ZN(_0468_)
);

AOI21_X1 _1585_ (
  .A(_0456_),
  .B1(_0468_),
  .B2(_0403_),
  .ZN(_0016_)
);

NOR2_X1 _1586_ (
  .A1(\ext_mult_res[17] ),
  .A2(_0373_),
  .ZN(_0469_)
);

INV_X1 _1587_ (
  .A(_1229_),
  .ZN(_0470_)
);

INV_X1 _1588_ (
  .A(_0467_),
  .ZN(_0471_)
);

NAND2_X1 _1589_ (
  .A1(_0451_),
  .A2(_0467_),
  .ZN(_0472_)
);

OAI221_X1 _1590_ (
  .A(_0470_),
  .B1(_0457_),
  .B2(_0471_),
  .C1(_0448_),
  .C2(_0472_),
  .ZN(_0473_)
);

INV_X1 _1591_ (
  .A(_0473_),
  .ZN(_0474_)
);

NOR2_X1 _1592_ (
  .A1(_0444_),
  .A2(_0472_),
  .ZN(_0475_)
);

NAND2_X1 _1593_ (
  .A1(_0429_),
  .A2(_0475_),
  .ZN(_0476_)
);

NAND3_X1 _1594_ (
  .A1(_0430_),
  .A2(_0475_),
  .A3(_0388_),
  .ZN(_0477_)
);

NAND3_X1 _1595_ (
  .A1(_0474_),
  .A2(_0476_),
  .A3(_0477_),
  .ZN(_0478_)
);

BUF_X1 _1596_ (
  .A(_1233_),
  .Z(_0479_)
);

XNOR2_X1 _1597_ (
  .A(_0478_),
  .B(_0479_),
  .ZN(_0480_)
);

AOI21_X1 _1598_ (
  .A(_0469_),
  .B1(_0480_),
  .B2(_0403_),
  .ZN(_0017_)
);

INV_X1 _1599_ (
  .A(_1061_),
  .ZN(_0481_)
);

INV_X1 _1600_ (
  .A(_1070_),
  .ZN(_0482_)
);

NAND2_X1 _1601_ (
  .A1(_0481_),
  .A2(_0482_),
  .ZN(_0483_)
);

NAND2_X1 _1602_ (
  .A1(_1061_),
  .A2(_1070_),
  .ZN(_0484_)
);

NAND2_X1 _1603_ (
  .A1(_0483_),
  .A2(_0484_),
  .ZN(_0485_)
);

INV_X1 _1604_ (
  .A(_0485_),
  .ZN(_0486_)
);

INV_X1 _1605_ (
  .A(_1081_),
  .ZN(_0487_)
);

NAND2_X1 _1606_ (
  .A1(_0487_),
  .A2(_1055_),
  .ZN(_0488_)
);

INV_X1 _1607_ (
  .A(_1055_),
  .ZN(_0489_)
);

NAND2_X1 _1608_ (
  .A1(_0489_),
  .A2(_1081_),
  .ZN(_0490_)
);

NAND2_X1 _1609_ (
  .A1(_0488_),
  .A2(_0490_),
  .ZN(_0491_)
);

NAND2_X1 _1610_ (
  .A1(_0486_),
  .A2(_0491_),
  .ZN(_0492_)
);

XNOR2_X1 _1611_ (
  .A(_1081_),
  .B(_1055_),
  .ZN(_0493_)
);

NAND2_X1 _1612_ (
  .A1(_0493_),
  .A2(_0485_),
  .ZN(_0494_)
);

NAND2_X1 _1613_ (
  .A1(_0492_),
  .A2(_0494_),
  .ZN(_0495_)
);

INV_X1 _1614_ (
  .A(_1224_),
  .ZN(_0496_)
);

NAND2_X1 _1615_ (
  .A1(_0496_),
  .A2(_1027_),
  .ZN(_0497_)
);

NAND2_X1 _1616_ (
  .A1(_1224_),
  .A2(_0987_),
  .ZN(_0498_)
);

XNOR2_X1 _1621_ (
  .A(_0495_),
  .B(_0502_),
  .ZN(_0503_)
);

INV_X1 _1622_ (
  .A(_1005_),
  .ZN(_0504_)
);

XNOR2_X1 _1623_ (
  .A(_0504_),
  .B(_1059_),
  .ZN(_0505_)
);

XNOR2_X1 _1624_ (
  .A(_1063_),
  .B(_1065_),
  .ZN(_0506_)
);

NAND2_X1 _1625_ (
  .A1(_0505_),
  .A2(_0506_),
  .ZN(_0507_)
);

NAND2_X1 _1626_ (
  .A1(_1063_),
  .A2(_1065_),
  .ZN(_0508_)
);

INV_X1 _1627_ (
  .A(_0508_),
  .ZN(_0509_)
);

NOR2_X1 _1628_ (
  .A1(_1063_),
  .A2(_1065_),
  .ZN(_0510_)
);

NOR2_X1 _1629_ (
  .A1(_0509_),
  .A2(_0510_),
  .ZN(_0511_)
);

XNOR2_X1 _1630_ (
  .A(_1005_),
  .B(_1059_),
  .ZN(_0512_)
);

NAND2_X1 _1631_ (
  .A1(_0511_),
  .A2(_0512_),
  .ZN(_0513_)
);

NAND2_X1 _1632_ (
  .A1(_0507_),
  .A2(_0513_),
  .ZN(_0514_)
);

INV_X1 _1633_ (
  .A(_0514_),
  .ZN(_0515_)
);

NAND2_X1 _1640_ (
  .A1(_0515_),
  .A2(_0521_),
  .ZN(_0522_)
);

NAND2_X1 _1645_ (
  .A1(_0526_),
  .A2(_0514_),
  .ZN(_0527_)
);

NAND2_X2 _1646_ (
  .A1(_0522_),
  .A2(_0527_),
  .ZN(_0528_)
);

NAND2_X1 _1647_ (
  .A1(_0503_),
  .A2(_0528_),
  .ZN(_0529_)
);

NAND2_X1 _1648_ (
  .A1(_0515_),
  .A2(_0526_),
  .ZN(_0530_)
);

NAND2_X1 _1649_ (
  .A1(_0521_),
  .A2(_0514_),
  .ZN(_0531_)
);

NAND2_X2 _1650_ (
  .A1(_0530_),
  .A2(_0531_),
  .ZN(_0532_)
);

XNOR2_X1 _1651_ (
  .A(_0491_),
  .B(_0485_),
  .ZN(_0533_)
);

NAND2_X1 _1652_ (
  .A1(_0533_),
  .A2(_0502_),
  .ZN(_0534_)
);

INV_X1 _1653_ (
  .A(_0502_),
  .ZN(_0535_)
);

NAND2_X1 _1654_ (
  .A1(_0495_),
  .A2(_0535_),
  .ZN(_0536_)
);

NAND2_X1 _1655_ (
  .A1(_0534_),
  .A2(_0536_),
  .ZN(_0537_)
);

NAND2_X1 _1656_ (
  .A1(_0532_),
  .A2(_0537_),
  .ZN(_0538_)
);

NAND2_X1 _1657_ (
  .A1(_0529_),
  .A2(_0538_),
  .ZN(_0539_)
);

OR2_X1 _1658_ (
  .A1(_1086_),
  .A2(_1078_),
  .ZN(_0540_)
);

NAND2_X1 _1659_ (
  .A1(_1078_),
  .A2(_1086_),
  .ZN(_0541_)
);

XOR2_X1 _1664_ (
  .A(_1068_),
  .B(_1231_),
  .Z(_0546_)
);

INV_X1 _1665_ (
  .A(_0546_),
  .ZN(_0547_)
);

NAND2_X2 _1666_ (
  .A1(_0545_),
  .A2(_0547_),
  .ZN(_0548_)
);

NAND2_X2 _1668_ (
  .A1(_0548_),
  .A2(_0549_),
  .ZN(_0550_)
);

XNOR2_X1 _1669_ (
  .A(_0967_),
  .B(_0903_),
  .ZN(_0551_)
);

XNOR2_X1 _1670_ (
  .A(_0874_),
  .B(_1073_),
  .ZN(_0552_)
);

XNOR2_X1 _1671_ (
  .A(_0551_),
  .B(_0552_),
  .ZN(_0553_)
);

INV_X1 _1672_ (
  .A(_0553_),
  .ZN(_0554_)
);

NAND2_X2 _1673_ (
  .A1(_0550_),
  .A2(_0554_),
  .ZN(_0555_)
);

NAND3_X1 _1674_ (
  .A1(_0548_),
  .A2(_0549_),
  .A3(_0553_),
  .ZN(_0556_)
);

NAND2_X2 _1675_ (
  .A1(_0555_),
  .A2(_0556_),
  .ZN(_0557_)
);

INV_X1 _1676_ (
  .A(_0557_),
  .ZN(_0558_)
);

NAND2_X2 _1677_ (
  .A1(_0539_),
  .A2(_0558_),
  .ZN(_0559_)
);

NAND2_X1 _1678_ (
  .A1(_0503_),
  .A2(_0532_),
  .ZN(_0560_)
);

NAND2_X1 _1679_ (
  .A1(_0528_),
  .A2(_0537_),
  .ZN(_0561_)
);

NAND2_X2 _1680_ (
  .A1(_0560_),
  .A2(_0561_),
  .ZN(_0562_)
);

NAND2_X2 _1681_ (
  .A1(_0562_),
  .A2(_0557_),
  .ZN(_0563_)
);

NAND2_X2 _1682_ (
  .A1(_0559_),
  .A2(_0563_),
  .ZN(_0564_)
);

INV_X1 _1683_ (
  .A(_0479_),
  .ZN(_0565_)
);

NOR3_X1 _1684_ (
  .A1(_0461_),
  .A2(_0471_),
  .A3(_0565_),
  .ZN(_0566_)
);

NAND3_X1 _1685_ (
  .A1(_0400_),
  .A2(_0440_),
  .A3(_0566_),
  .ZN(_0567_)
);

NAND3_X1 _1686_ (
  .A1(_0459_),
  .A2(_0467_),
  .A3(_0479_),
  .ZN(_0568_)
);

INV_X1 _1687_ (
  .A(_1232_),
  .ZN(_0569_)
);

NAND2_X1 _1688_ (
  .A1(_0479_),
  .A2(_1229_),
  .ZN(_0570_)
);

NAND3_X1 _1689_ (
  .A1(_0568_),
  .A2(_0569_),
  .A3(_0570_),
  .ZN(_0571_)
);

INV_X1 _1690_ (
  .A(_0571_),
  .ZN(_0572_)
);

NAND2_X1 _1691_ (
  .A1(_0439_),
  .A2(_0566_),
  .ZN(_0573_)
);

AND3_X1 _1692_ (
  .A1(_0567_),
  .A2(_0572_),
  .A3(_0573_),
  .ZN(_0574_)
);

INV_X1 _1693_ (
  .A(_0574_),
  .ZN(_0575_)
);

NAND2_X2 _1694_ (
  .A1(_0564_),
  .A2(_0575_),
  .ZN(_0576_)
);

NAND3_X1 _1695_ (
  .A1(_0559_),
  .A2(_0563_),
  .A3(_0574_),
  .ZN(_0577_)
);

NAND3_X1 _1696_ (
  .A1(_0576_),
  .A2(_0577_),
  .A3(_0374_),
  .ZN(_0578_)
);

NAND2_X1 _1697_ (
  .A1(_0387_),
  .A2(\ext_mult_res[18] ),
  .ZN(_0579_)
);

NAND2_X1 _1698_ (
  .A1(_0578_),
  .A2(_0579_),
  .ZN(_0018_)
);

NAND2_X1 _1699_ (
  .A1(_0385_),
  .A2(result[0]),
  .ZN(_0580_)
);

BUF_X1 _1700_ (
  .A(dclr),
  .Z(_0581_)
);

OAI21_X1 _1701_ (
  .A(_0368_),
  .B1(_1089_),
  .B2(_0581_),
  .ZN(_0582_)
);

INV_X1 _1702_ (
  .A(_0581_),
  .ZN(_0583_)
);

BUF_X1 _1703_ (
  .A(_0583_),
  .Z(_0584_)
);

NOR2_X1 _1704_ (
  .A1(_0584_),
  .A2(\ext_mult_res[0] ),
  .ZN(_0585_)
);

OAI21_X1 _1705_ (
  .A(_0580_),
  .B1(_0582_),
  .B2(_0585_),
  .ZN(_0019_)
);

NAND2_X1 _1706_ (
  .A1(_0385_),
  .A2(result[1]),
  .ZN(_0586_)
);

OAI21_X1 _1707_ (
  .A(_0368_),
  .B1(_0581_),
  .B2(_0680_),
  .ZN(_0587_)
);

NOR2_X1 _1708_ (
  .A1(_0584_),
  .A2(\ext_mult_res[1] ),
  .ZN(_0588_)
);

OAI21_X1 _1709_ (
  .A(_0586_),
  .B1(_0587_),
  .B2(_0588_),
  .ZN(_0020_)
);

INV_X1 _1710_ (
  .A(_1093_),
  .ZN(_0589_)
);

NOR2_X1 _1711_ (
  .A1(_0589_),
  .A2(_0679_),
  .ZN(_0590_)
);

INV_X1 _1712_ (
  .A(_0590_),
  .ZN(_0591_)
);

NAND2_X1 _1713_ (
  .A1(_0589_),
  .A2(_0679_),
  .ZN(_0592_)
);

NAND3_X1 _1714_ (
  .A1(_0591_),
  .A2(_0583_),
  .A3(_0592_),
  .ZN(_0593_)
);

BUF_X2 _1715_ (
  .A(_0583_),
  .Z(_0594_)
);

OAI21_X1 _1716_ (
  .A(_0593_),
  .B1(_0594_),
  .B2(_0376_),
  .ZN(_0595_)
);

MUX2_X1 _1717_ (
  .A(result[2]),
  .B(_0595_),
  .S(_0373_),
  .Z(_0021_)
);

OAI21_X1 _1718_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(_0378_),
  .ZN(_0596_)
);

NAND2_X1 _1719_ (
  .A1(_1088_),
  .A2(_1091_),
  .ZN(_0597_)
);

INV_X1 _1720_ (
  .A(_1090_),
  .ZN(_0598_)
);

INV_X1 _1721_ (
  .A(_1092_),
  .ZN(_0599_)
);

NAND3_X1 _1722_ (
  .A1(_0597_),
  .A2(_0598_),
  .A3(_0599_),
  .ZN(_0600_)
);

NAND2_X1 _1723_ (
  .A1(_0589_),
  .A2(_0599_),
  .ZN(_0601_)
);

NAND2_X1 _1724_ (
  .A1(_0600_),
  .A2(_0601_),
  .ZN(_0602_)
);

XNOR2_X1 _1725_ (
  .A(_0602_),
  .B(_1095_),
  .ZN(_0603_)
);

BUF_X1 _1726_ (
  .A(_0583_),
  .Z(_0604_)
);

AOI21_X1 _1727_ (
  .A(_0596_),
  .B1(_0603_),
  .B2(_0604_),
  .ZN(_0605_)
);

INV_X1 _1728_ (
  .A(result[3]),
  .ZN(_0606_)
);

AOI21_X1 _1729_ (
  .A(_0605_),
  .B1(_0606_),
  .B2(_0387_),
  .ZN(_0022_)
);

OAI21_X1 _1730_ (
  .A(_0367_),
  .B1(_0583_),
  .B2(_0380_),
  .ZN(_0607_)
);

INV_X1 _1731_ (
  .A(_1094_),
  .ZN(_0608_)
);

INV_X1 _1732_ (
  .A(_1095_),
  .ZN(_0609_)
);

OAI21_X1 _1733_ (
  .A(_0608_),
  .B1(_0609_),
  .B2(_0599_),
  .ZN(_0610_)
);

INV_X1 _1734_ (
  .A(_0610_),
  .ZN(_0611_)
);

OAI21_X4 _1735_ (
  .A(_0611_),
  .B1(_0609_),
  .B2(_0591_),
  .ZN(_0612_)
);

INV_X1 _1736_ (
  .A(_1097_),
  .ZN(_0613_)
);

XNOR2_X1 _1737_ (
  .A(_0612_),
  .B(_0613_),
  .ZN(_0614_)
);

AOI21_X1 _1738_ (
  .A(_0607_),
  .B1(_0614_),
  .B2(_0604_),
  .ZN(_0615_)
);

INV_X1 _1739_ (
  .A(result[4]),
  .ZN(_0616_)
);

AOI21_X1 _1740_ (
  .A(_0615_),
  .B1(_0616_),
  .B2(_0387_),
  .ZN(_0023_)
);

NAND2_X1 _1741_ (
  .A1(_1095_),
  .A2(_1097_),
  .ZN(_0617_)
);

INV_X1 _1742_ (
  .A(_0617_),
  .ZN(_0618_)
);

NAND3_X1 _1743_ (
  .A1(_0600_),
  .A2(_0601_),
  .A3(_0618_),
  .ZN(_0619_)
);

INV_X1 _1744_ (
  .A(_1096_),
  .ZN(_0620_)
);

OAI21_X1 _1745_ (
  .A(_0620_),
  .B1(_0613_),
  .B2(_0608_),
  .ZN(_0621_)
);

INV_X1 _1746_ (
  .A(_0621_),
  .ZN(_0622_)
);

NAND2_X1 _1747_ (
  .A1(_0619_),
  .A2(_0622_),
  .ZN(_0623_)
);

BUF_X2 _1748_ (
  .A(_1099_),
  .Z(_0624_)
);

XNOR2_X1 _1749_ (
  .A(_0623_),
  .B(_0624_),
  .ZN(_0625_)
);

AOI21_X1 _1750_ (
  .A(_0385_),
  .B1(_0625_),
  .B2(_0594_),
  .ZN(_0626_)
);

OAI21_X1 _1751_ (
  .A(_0626_),
  .B1(_0584_),
  .B2(\ext_mult_res[5] ),
  .ZN(_0627_)
);

INV_X1 _1752_ (
  .A(result[5]),
  .ZN(_0628_)
);

OAI21_X1 _1753_ (
  .A(_0627_),
  .B1(_0403_),
  .B2(_0628_),
  .ZN(_0024_)
);

INV_X1 _1754_ (
  .A(_1098_),
  .ZN(_0629_)
);

INV_X1 _1755_ (
  .A(_0624_),
  .ZN(_0630_)
);

OAI21_X1 _1756_ (
  .A(_0629_),
  .B1(_0630_),
  .B2(_0620_),
  .ZN(_0631_)
);

INV_X1 _1757_ (
  .A(_0631_),
  .ZN(_0632_)
);

INV_X1 _1758_ (
  .A(_0612_),
  .ZN(_0633_)
);

NAND2_X1 _1759_ (
  .A1(_1097_),
  .A2(_0624_),
  .ZN(_0634_)
);

OAI21_X1 _1760_ (
  .A(_0632_),
  .B1(_0633_),
  .B2(_0634_),
  .ZN(_0635_)
);

CLKBUF_X2 _1761_ (
  .A(_1101_),
  .Z(_0636_)
);

XNOR2_X1 _1762_ (
  .A(_0635_),
  .B(_0636_),
  .ZN(_0041_)
);

NAND2_X1 _1763_ (
  .A1(_0041_),
  .A2(_0604_),
  .ZN(_0042_)
);

NAND2_X1 _1764_ (
  .A1(_0382_),
  .A2(_0581_),
  .ZN(_0043_)
);

NAND3_X1 _1765_ (
  .A1(_0042_),
  .A2(_0374_),
  .A3(_0043_),
  .ZN(_0044_)
);

INV_X1 _1766_ (
  .A(result[6]),
  .ZN(_0045_)
);

OAI21_X1 _1767_ (
  .A(_0044_),
  .B1(_0403_),
  .B2(_0045_),
  .ZN(_0025_)
);

NAND2_X1 _1768_ (
  .A1(_0636_),
  .A2(_1098_),
  .ZN(_0046_)
);

INV_X1 _1769_ (
  .A(_1100_),
  .ZN(_0047_)
);

NAND2_X1 _1770_ (
  .A1(_0046_),
  .A2(_0047_),
  .ZN(_0048_)
);

INV_X1 _1771_ (
  .A(_0048_),
  .ZN(_0049_)
);

NAND2_X1 _1772_ (
  .A1(_0624_),
  .A2(_0636_),
  .ZN(_0050_)
);

OAI21_X1 _1773_ (
  .A(_0049_),
  .B1(_0622_),
  .B2(_0050_),
  .ZN(_0051_)
);

INV_X1 _1774_ (
  .A(_0051_),
  .ZN(_0052_)
);

OAI21_X1 _1775_ (
  .A(_0052_),
  .B1(_0619_),
  .B2(_0050_),
  .ZN(_0053_)
);

BUF_X2 _1776_ (
  .A(_1103_),
  .Z(_0054_)
);

XNOR2_X1 _1777_ (
  .A(_0053_),
  .B(_0054_),
  .ZN(_0055_)
);

NAND2_X1 _1778_ (
  .A1(_0055_),
  .A2(_0604_),
  .ZN(_0056_)
);

NAND2_X1 _1779_ (
  .A1(_0384_),
  .A2(_0581_),
  .ZN(_0057_)
);

NAND3_X1 _1780_ (
  .A1(_0056_),
  .A2(_0374_),
  .A3(_0057_),
  .ZN(_0058_)
);

INV_X1 _1781_ (
  .A(result[7]),
  .ZN(_0059_)
);

OAI21_X1 _1782_ (
  .A(_0058_),
  .B1(_0403_),
  .B2(_0059_),
  .ZN(_0026_)
);

NAND2_X1 _1783_ (
  .A1(_0385_),
  .A2(result[8]),
  .ZN(_0060_)
);

INV_X1 _1784_ (
  .A(_1102_),
  .ZN(_0061_)
);

INV_X1 _1785_ (
  .A(_0054_),
  .ZN(_0062_)
);

OAI21_X1 _1786_ (
  .A(_0061_),
  .B1(_0062_),
  .B2(_0047_),
  .ZN(_0063_)
);

INV_X1 _1787_ (
  .A(_0063_),
  .ZN(_0064_)
);

NAND2_X1 _1788_ (
  .A1(_0636_),
  .A2(_0054_),
  .ZN(_0065_)
);

OAI21_X1 _1789_ (
  .A(_0064_),
  .B1(_0632_),
  .B2(_0065_),
  .ZN(_0066_)
);

INV_X1 _1790_ (
  .A(_0066_),
  .ZN(_0067_)
);

NOR2_X1 _1791_ (
  .A1(_0634_),
  .A2(_0065_),
  .ZN(_0068_)
);

INV_X1 _1792_ (
  .A(_0068_),
  .ZN(_0069_)
);

OAI21_X1 _1793_ (
  .A(_0067_),
  .B1(_0633_),
  .B2(_0069_),
  .ZN(_0070_)
);

INV_X1 _1794_ (
  .A(_1105_),
  .ZN(_0071_)
);

XNOR2_X1 _1795_ (
  .A(_0070_),
  .B(_0071_),
  .ZN(_0072_)
);

OAI21_X1 _1796_ (
  .A(_0368_),
  .B1(_0072_),
  .B2(_0581_),
  .ZN(_0073_)
);

NOR2_X1 _1797_ (
  .A1(_0584_),
  .A2(\ext_mult_res[8] ),
  .ZN(_0074_)
);

OAI21_X1 _1798_ (
  .A(_0060_),
  .B1(_0073_),
  .B2(_0074_),
  .ZN(_0027_)
);

OAI21_X1 _1799_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[9] ),
  .ZN(_0075_)
);

INV_X1 _1800_ (
  .A(_0075_),
  .ZN(_0076_)
);

NAND2_X2 _1801_ (
  .A1(_0054_),
  .A2(_1105_),
  .ZN(_0077_)
);

INV_X1 _1802_ (
  .A(_0077_),
  .ZN(_0078_)
);

NAND2_X1 _1803_ (
  .A1(_0053_),
  .A2(_0078_),
  .ZN(_0079_)
);

INV_X1 _1804_ (
  .A(_1104_),
  .ZN(_0080_)
);

OAI21_X1 _1805_ (
  .A(_0080_),
  .B1(_0071_),
  .B2(_0061_),
  .ZN(_0081_)
);

INV_X1 _1806_ (
  .A(_0081_),
  .ZN(_0082_)
);

NAND2_X1 _1807_ (
  .A1(_0079_),
  .A2(_0082_),
  .ZN(_0083_)
);

INV_X1 _1808_ (
  .A(_1107_),
  .ZN(_0084_)
);

XNOR2_X1 _1809_ (
  .A(_0083_),
  .B(_0084_),
  .ZN(_0085_)
);

OAI21_X1 _1810_ (
  .A(_0076_),
  .B1(_0085_),
  .B2(_0581_),
  .ZN(_0086_)
);

NAND2_X1 _1811_ (
  .A1(_0387_),
  .A2(result[9]),
  .ZN(_0087_)
);

NAND2_X1 _1812_ (
  .A1(_0086_),
  .A2(_0087_),
  .ZN(_0028_)
);

NAND2_X1 _1813_ (
  .A1(_0385_),
  .A2(result[10]),
  .ZN(_0088_)
);

OAI21_X1 _1814_ (
  .A(_0632_),
  .B1(_0611_),
  .B2(_0634_),
  .ZN(_0089_)
);

NAND2_X1 _1815_ (
  .A1(_1105_),
  .A2(_1107_),
  .ZN(_0090_)
);

NOR2_X1 _1816_ (
  .A1(_0065_),
  .A2(_0090_),
  .ZN(_0091_)
);

NAND2_X1 _1817_ (
  .A1(_0089_),
  .A2(_0091_),
  .ZN(_0092_)
);

INV_X1 _1818_ (
  .A(_1106_),
  .ZN(_0093_)
);

OAI21_X1 _1819_ (
  .A(_0093_),
  .B1(_0084_),
  .B2(_0080_),
  .ZN(_0094_)
);

INV_X1 _1820_ (
  .A(_0094_),
  .ZN(_0095_)
);

OAI21_X1 _1821_ (
  .A(_0095_),
  .B1(_0064_),
  .B2(_0090_),
  .ZN(_0096_)
);

INV_X1 _1822_ (
  .A(_0096_),
  .ZN(_0097_)
);

NOR3_X1 _1823_ (
  .A1(_0634_),
  .A2(_0589_),
  .A3(_0609_),
  .ZN(_0098_)
);

INV_X1 _1824_ (
  .A(_0679_),
  .ZN(_0099_)
);

NAND3_X1 _1825_ (
  .A1(_0098_),
  .A2(_0099_),
  .A3(_0091_),
  .ZN(_0100_)
);

NAND3_X1 _1826_ (
  .A1(_0092_),
  .A2(_0097_),
  .A3(_0100_),
  .ZN(_0101_)
);

INV_X1 _1827_ (
  .A(_1109_),
  .ZN(_0102_)
);

XNOR2_X1 _1828_ (
  .A(_0101_),
  .B(_0102_),
  .ZN(_0103_)
);

NOR2_X1 _1829_ (
  .A1(_0103_),
  .A2(_0581_),
  .ZN(_0104_)
);

OAI21_X1 _1830_ (
  .A(_0368_),
  .B1(_0584_),
  .B2(\ext_mult_res[10] ),
  .ZN(_0105_)
);

OAI21_X1 _1831_ (
  .A(_0088_),
  .B1(_0104_),
  .B2(_0105_),
  .ZN(_0029_)
);

NAND2_X1 _1832_ (
  .A1(_0385_),
  .A2(result[11]),
  .ZN(_0106_)
);

NAND2_X1 _1833_ (
  .A1(_1107_),
  .A2(_1109_),
  .ZN(_0107_)
);

NOR2_X2 _1834_ (
  .A1(_0077_),
  .A2(_0107_),
  .ZN(_0108_)
);

NAND2_X1 _1835_ (
  .A1(_0051_),
  .A2(_0108_),
  .ZN(_0109_)
);

INV_X1 _1836_ (
  .A(_1108_),
  .ZN(_0110_)
);

OAI21_X1 _1837_ (
  .A(_0110_),
  .B1(_0102_),
  .B2(_0093_),
  .ZN(_0111_)
);

INV_X1 _1838_ (
  .A(_0111_),
  .ZN(_0112_)
);

OAI21_X1 _1839_ (
  .A(_0112_),
  .B1(_0082_),
  .B2(_0107_),
  .ZN(_0113_)
);

INV_X1 _1840_ (
  .A(_0113_),
  .ZN(_0114_)
);

NAND2_X1 _1841_ (
  .A1(_0109_),
  .A2(_0114_),
  .ZN(_0115_)
);

INV_X1 _1842_ (
  .A(_0115_),
  .ZN(_0116_)
);

NAND4_X1 _1843_ (
  .A1(_0108_),
  .A2(_0618_),
  .A3(_0636_),
  .A4(_0624_),
  .ZN(_0117_)
);

INV_X1 _1844_ (
  .A(_0117_),
  .ZN(_0118_)
);

INV_X1 _1845_ (
  .A(_0602_),
  .ZN(_0119_)
);

NAND2_X1 _1846_ (
  .A1(_0118_),
  .A2(_0119_),
  .ZN(_0120_)
);

NAND2_X1 _1847_ (
  .A1(_0116_),
  .A2(_0120_),
  .ZN(_0121_)
);

INV_X1 _1848_ (
  .A(_1111_),
  .ZN(_0122_)
);

NAND2_X1 _1849_ (
  .A1(_0121_),
  .A2(_0122_),
  .ZN(_0123_)
);

NAND3_X1 _1850_ (
  .A1(_0116_),
  .A2(_1111_),
  .A3(_0120_),
  .ZN(_0124_)
);

NAND3_X1 _1851_ (
  .A1(_0123_),
  .A2(_0124_),
  .A3(_0604_),
  .ZN(_0125_)
);

NAND2_X1 _1852_ (
  .A1(_0125_),
  .A2(_0374_),
  .ZN(_0126_)
);

NOR2_X1 _1853_ (
  .A1(_0584_),
  .A2(\ext_mult_res[11] ),
  .ZN(_0127_)
);

OAI21_X1 _1854_ (
  .A(_0106_),
  .B1(_0126_),
  .B2(_0127_),
  .ZN(_0030_)
);

NAND2_X1 _1855_ (
  .A1(_0385_),
  .A2(result[12]),
  .ZN(_0128_)
);

NAND2_X1 _1856_ (
  .A1(_1109_),
  .A2(_1111_),
  .ZN(_0129_)
);

NOR2_X1 _1857_ (
  .A1(_0090_),
  .A2(_0129_),
  .ZN(_0130_)
);

NAND2_X1 _1858_ (
  .A1(_0066_),
  .A2(_0130_),
  .ZN(_0131_)
);

INV_X1 _1859_ (
  .A(_1110_),
  .ZN(_0132_)
);

OAI21_X1 _1860_ (
  .A(_0132_),
  .B1(_0122_),
  .B2(_0110_),
  .ZN(_0133_)
);

INV_X1 _1861_ (
  .A(_0133_),
  .ZN(_0134_)
);

OAI21_X1 _1862_ (
  .A(_0134_),
  .B1(_0095_),
  .B2(_0129_),
  .ZN(_0135_)
);

INV_X1 _1863_ (
  .A(_0135_),
  .ZN(_0136_)
);

NAND2_X1 _1864_ (
  .A1(_0131_),
  .A2(_0136_),
  .ZN(_0137_)
);

INV_X1 _1865_ (
  .A(_0137_),
  .ZN(_0138_)
);

NAND2_X1 _1866_ (
  .A1(_0068_),
  .A2(_0130_),
  .ZN(_0139_)
);

INV_X1 _1867_ (
  .A(_0139_),
  .ZN(_0140_)
);

NAND2_X1 _1868_ (
  .A1(_0612_),
  .A2(_0140_),
  .ZN(_0141_)
);

NAND2_X1 _1869_ (
  .A1(_0138_),
  .A2(_0141_),
  .ZN(_0142_)
);

INV_X1 _1870_ (
  .A(_1113_),
  .ZN(_0143_)
);

NAND2_X1 _1871_ (
  .A1(_0142_),
  .A2(_0143_),
  .ZN(_0144_)
);

NAND3_X1 _1872_ (
  .A1(_0138_),
  .A2(_1113_),
  .A3(_0141_),
  .ZN(_0145_)
);

AND3_X1 _1873_ (
  .A1(_0144_),
  .A2(_0145_),
  .A3(_0594_),
  .ZN(_0146_)
);

OAI21_X1 _1874_ (
  .A(_0368_),
  .B1(_0584_),
  .B2(\ext_mult_res[12] ),
  .ZN(_0147_)
);

OAI21_X1 _1875_ (
  .A(_0128_),
  .B1(_0146_),
  .B2(_0147_),
  .ZN(_0031_)
);

NAND2_X1 _1876_ (
  .A1(_0385_),
  .A2(result[13]),
  .ZN(_0148_)
);

NAND2_X1 _1877_ (
  .A1(_0048_),
  .A2(_0078_),
  .ZN(_0149_)
);

NAND2_X1 _1878_ (
  .A1(_0082_),
  .A2(_0149_),
  .ZN(_0150_)
);

NAND2_X1 _1879_ (
  .A1(_1111_),
  .A2(_1113_),
  .ZN(_0151_)
);

NOR2_X1 _1880_ (
  .A1(_0107_),
  .A2(_0151_),
  .ZN(_0152_)
);

NAND2_X1 _1881_ (
  .A1(_0150_),
  .A2(_0152_),
  .ZN(_0153_)
);

INV_X1 _1882_ (
  .A(_0151_),
  .ZN(_0154_)
);

NAND2_X1 _1883_ (
  .A1(_0111_),
  .A2(_0154_),
  .ZN(_0155_)
);

INV_X1 _1884_ (
  .A(_1112_),
  .ZN(_0156_)
);

OAI21_X1 _1885_ (
  .A(_0156_),
  .B1(_0143_),
  .B2(_0132_),
  .ZN(_0157_)
);

INV_X1 _1886_ (
  .A(_0157_),
  .ZN(_0158_)
);

NAND2_X1 _1887_ (
  .A1(_0155_),
  .A2(_0158_),
  .ZN(_0159_)
);

INV_X1 _1888_ (
  .A(_0159_),
  .ZN(_0160_)
);

NAND2_X1 _1889_ (
  .A1(_0153_),
  .A2(_0160_),
  .ZN(_0161_)
);

INV_X1 _1890_ (
  .A(_0161_),
  .ZN(_0162_)
);

INV_X1 _1891_ (
  .A(_0623_),
  .ZN(_0163_)
);

NOR2_X2 _1892_ (
  .A1(_0050_),
  .A2(_0077_),
  .ZN(_0164_)
);

NAND2_X1 _1893_ (
  .A1(_0164_),
  .A2(_0152_),
  .ZN(_0165_)
);

OAI21_X1 _1894_ (
  .A(_0162_),
  .B1(_0163_),
  .B2(_0165_),
  .ZN(_0166_)
);

INV_X1 _1895_ (
  .A(_1115_),
  .ZN(_0167_)
);

XNOR2_X1 _1896_ (
  .A(_0166_),
  .B(_0167_),
  .ZN(_0168_)
);

NOR2_X1 _1897_ (
  .A1(_0168_),
  .A2(_0581_),
  .ZN(_0169_)
);

OAI21_X1 _1898_ (
  .A(_0368_),
  .B1(_0604_),
  .B2(\ext_mult_res[13] ),
  .ZN(_0170_)
);

OAI21_X1 _1899_ (
  .A(_0148_),
  .B1(_0169_),
  .B2(_0170_),
  .ZN(_0032_)
);

NAND2_X1 _1900_ (
  .A1(_1113_),
  .A2(_1115_),
  .ZN(_0171_)
);

NOR2_X1 _1901_ (
  .A1(_0129_),
  .A2(_0171_),
  .ZN(_0172_)
);

NAND3_X1 _1902_ (
  .A1(_0635_),
  .A2(_0091_),
  .A3(_0172_),
  .ZN(_0173_)
);

INV_X1 _1903_ (
  .A(_1114_),
  .ZN(_0174_)
);

OAI21_X1 _1904_ (
  .A(_0174_),
  .B1(_0167_),
  .B2(_0156_),
  .ZN(_0175_)
);

INV_X1 _1905_ (
  .A(_0175_),
  .ZN(_0176_)
);

OAI21_X1 _1906_ (
  .A(_0176_),
  .B1(_0134_),
  .B2(_0171_),
  .ZN(_0177_)
);

AOI21_X1 _1907_ (
  .A(_0177_),
  .B1(_0172_),
  .B2(_0096_),
  .ZN(_0178_)
);

NAND2_X1 _1908_ (
  .A1(_0173_),
  .A2(_0178_),
  .ZN(_0179_)
);

INV_X1 _1909_ (
  .A(_1117_),
  .ZN(_0180_)
);

NAND2_X1 _1910_ (
  .A1(_0179_),
  .A2(_0180_),
  .ZN(_0181_)
);

NAND3_X1 _1911_ (
  .A1(_0173_),
  .A2(_1117_),
  .A3(_0178_),
  .ZN(_0182_)
);

NAND3_X1 _1912_ (
  .A1(_0181_),
  .A2(_0182_),
  .A3(_0604_),
  .ZN(_0183_)
);

OAI21_X1 _1913_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[14] ),
  .ZN(_0184_)
);

INV_X1 _1914_ (
  .A(_0184_),
  .ZN(_0185_)
);

NAND2_X1 _1915_ (
  .A1(_0183_),
  .A2(_0185_),
  .ZN(_0186_)
);

NAND2_X1 _1916_ (
  .A1(_0387_),
  .A2(result[14]),
  .ZN(_0187_)
);

NAND2_X1 _1917_ (
  .A1(_0186_),
  .A2(_0187_),
  .ZN(_0033_)
);

NAND2_X1 _1918_ (
  .A1(_1115_),
  .A2(_1117_),
  .ZN(_0188_)
);

NOR2_X1 _1919_ (
  .A1(_0151_),
  .A2(_0188_),
  .ZN(_0189_)
);

NAND3_X1 _1920_ (
  .A1(_0053_),
  .A2(_0108_),
  .A3(_0189_),
  .ZN(_0190_)
);

INV_X1 _1921_ (
  .A(_1116_),
  .ZN(_0191_)
);

OAI21_X1 _1922_ (
  .A(_0191_),
  .B1(_0180_),
  .B2(_0174_),
  .ZN(_0192_)
);

INV_X1 _1923_ (
  .A(_0192_),
  .ZN(_0193_)
);

OAI21_X1 _1924_ (
  .A(_0193_),
  .B1(_0158_),
  .B2(_0188_),
  .ZN(_0194_)
);

AOI21_X1 _1925_ (
  .A(_0194_),
  .B1(_0189_),
  .B2(_0113_),
  .ZN(_0195_)
);

NAND2_X1 _1926_ (
  .A1(_0190_),
  .A2(_0195_),
  .ZN(_0196_)
);

INV_X1 _1927_ (
  .A(_1119_),
  .ZN(_0197_)
);

NAND2_X1 _1928_ (
  .A1(_0196_),
  .A2(_0197_),
  .ZN(_0198_)
);

NAND3_X1 _1929_ (
  .A1(_0190_),
  .A2(_1119_),
  .A3(_0195_),
  .ZN(_0199_)
);

NAND3_X1 _1930_ (
  .A1(_0198_),
  .A2(_0199_),
  .A3(_0604_),
  .ZN(_0200_)
);

OAI21_X1 _1931_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[15] ),
  .ZN(_0201_)
);

INV_X1 _1932_ (
  .A(_0201_),
  .ZN(_0202_)
);

NAND2_X1 _1933_ (
  .A1(_0200_),
  .A2(_0202_),
  .ZN(_0203_)
);

NAND2_X1 _1934_ (
  .A1(_0387_),
  .A2(result[15]),
  .ZN(_0204_)
);

NAND2_X1 _1935_ (
  .A1(_0203_),
  .A2(_0204_),
  .ZN(_0034_)
);

OAI21_X1 _1936_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[16] ),
  .ZN(_0205_)
);

INV_X1 _1937_ (
  .A(_0205_),
  .ZN(_0206_)
);

NAND2_X1 _1938_ (
  .A1(_1117_),
  .A2(_1119_),
  .ZN(_0207_)
);

NOR2_X1 _1939_ (
  .A1(_0171_),
  .A2(_0207_),
  .ZN(_0208_)
);

NAND3_X1 _1940_ (
  .A1(_0070_),
  .A2(_0130_),
  .A3(_0208_),
  .ZN(_0209_)
);

BUF_X2 _1941_ (
  .A(_1121_),
  .Z(_0210_)
);

INV_X1 _1942_ (
  .A(_1118_),
  .ZN(_0211_)
);

OAI21_X1 _1943_ (
  .A(_0211_),
  .B1(_0197_),
  .B2(_0191_),
  .ZN(_0212_)
);

INV_X1 _1944_ (
  .A(_0212_),
  .ZN(_0213_)
);

OAI21_X1 _1945_ (
  .A(_0213_),
  .B1(_0176_),
  .B2(_0207_),
  .ZN(_0214_)
);

AOI21_X1 _1946_ (
  .A(_0214_),
  .B1(_0208_),
  .B2(_0135_),
  .ZN(_0215_)
);

NAND3_X1 _1947_ (
  .A1(_0209_),
  .A2(_0210_),
  .A3(_0215_),
  .ZN(_0216_)
);

NAND2_X1 _1948_ (
  .A1(_0216_),
  .A2(_0604_),
  .ZN(_0217_)
);

AOI21_X1 _1949_ (
  .A(_0210_),
  .B1(_0209_),
  .B2(_0215_),
  .ZN(_0218_)
);

OAI21_X1 _1950_ (
  .A(_0206_),
  .B1(_0217_),
  .B2(_0218_),
  .ZN(_0219_)
);

NAND2_X1 _1951_ (
  .A1(_0387_),
  .A2(result[16]),
  .ZN(_0220_)
);

NAND2_X1 _1952_ (
  .A1(_0219_),
  .A2(_0220_),
  .ZN(_0035_)
);

OAI21_X1 _1953_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[17] ),
  .ZN(_0221_)
);

INV_X1 _1954_ (
  .A(_0221_),
  .ZN(_0222_)
);

OAI21_X1 _1955_ (
  .A(_0599_),
  .B1(_0589_),
  .B2(_0598_),
  .ZN(_0223_)
);

INV_X1 _1956_ (
  .A(_0223_),
  .ZN(_0224_)
);

OAI21_X1 _1957_ (
  .A(_0622_),
  .B1(_0224_),
  .B2(_0617_),
  .ZN(_0225_)
);

NAND2_X1 _1958_ (
  .A1(_0225_),
  .A2(_0164_),
  .ZN(_0226_)
);

INV_X1 _1959_ (
  .A(_0150_),
  .ZN(_0227_)
);

NAND2_X1 _1960_ (
  .A1(_0226_),
  .A2(_0227_),
  .ZN(_0228_)
);

NAND2_X2 _1961_ (
  .A1(_1119_),
  .A2(_0210_),
  .ZN(_0229_)
);

NOR2_X2 _1962_ (
  .A1(_0188_),
  .A2(_0229_),
  .ZN(_0230_)
);

AND2_X1 _1963_ (
  .A1(_0152_),
  .A2(_0230_),
  .ZN(_0231_)
);

NAND2_X1 _1964_ (
  .A1(_0228_),
  .A2(_0231_),
  .ZN(_0232_)
);

INV_X1 _1965_ (
  .A(_0229_),
  .ZN(_0233_)
);

NAND2_X1 _1966_ (
  .A1(_0192_),
  .A2(_0233_),
  .ZN(_0234_)
);

INV_X1 _1967_ (
  .A(_1120_),
  .ZN(_0235_)
);

INV_X1 _1968_ (
  .A(_0210_),
  .ZN(_0236_)
);

OAI21_X1 _1969_ (
  .A(_0235_),
  .B1(_0236_),
  .B2(_0211_),
  .ZN(_0237_)
);

INV_X1 _1970_ (
  .A(_0237_),
  .ZN(_0238_)
);

NAND2_X1 _1971_ (
  .A1(_0234_),
  .A2(_0238_),
  .ZN(_0239_)
);

AOI21_X1 _1972_ (
  .A(_0239_),
  .B1(_0230_),
  .B2(_0159_),
  .ZN(_0240_)
);

AND3_X1 _1973_ (
  .A1(_0618_),
  .A2(_1091_),
  .A3(_1093_),
  .ZN(_0241_)
);

NAND4_X1 _1974_ (
  .A1(_0231_),
  .A2(_0241_),
  .A3(_0164_),
  .A4(_1088_),
  .ZN(_0242_)
);

NAND3_X1 _1975_ (
  .A1(_0232_),
  .A2(_0240_),
  .A3(_0242_),
  .ZN(_0243_)
);

INV_X1 _1976_ (
  .A(_1123_),
  .ZN(_0244_)
);

NAND2_X1 _1977_ (
  .A1(_0243_),
  .A2(_0244_),
  .ZN(_0245_)
);

NAND2_X1 _1978_ (
  .A1(_0245_),
  .A2(_0604_),
  .ZN(_0246_)
);

NOR2_X1 _1979_ (
  .A1(_0243_),
  .A2(_0244_),
  .ZN(_0247_)
);

OAI21_X1 _1980_ (
  .A(_0222_),
  .B1(_0246_),
  .B2(_0247_),
  .ZN(_0248_)
);

NAND2_X1 _1981_ (
  .A1(_0387_),
  .A2(result[17]),
  .ZN(_0249_)
);

NAND2_X1 _1982_ (
  .A1(_0248_),
  .A2(_0249_),
  .ZN(_0036_)
);

NOR2_X1 _1983_ (
  .A1(_0368_),
  .A2(result[18]),
  .ZN(_0250_)
);

NAND2_X1 _1984_ (
  .A1(_0092_),
  .A2(_0097_),
  .ZN(_0251_)
);

NAND2_X1 _1985_ (
  .A1(_0210_),
  .A2(_1123_),
  .ZN(_0252_)
);

NOR2_X1 _1986_ (
  .A1(_0207_),
  .A2(_0252_),
  .ZN(_0253_)
);

AND2_X1 _1987_ (
  .A1(_0172_),
  .A2(_0253_),
  .ZN(_0254_)
);

NAND2_X1 _1988_ (
  .A1(_0251_),
  .A2(_0254_),
  .ZN(_0255_)
);

INV_X1 _1989_ (
  .A(_1122_),
  .ZN(_0256_)
);

OAI21_X1 _1990_ (
  .A(_0256_),
  .B1(_0244_),
  .B2(_0235_),
  .ZN(_0257_)
);

INV_X1 _1991_ (
  .A(_0257_),
  .ZN(_0258_)
);

OAI21_X1 _1992_ (
  .A(_0258_),
  .B1(_0213_),
  .B2(_0252_),
  .ZN(_0259_)
);

AOI21_X1 _1993_ (
  .A(_0259_),
  .B1(_0253_),
  .B2(_0177_),
  .ZN(_0260_)
);

NAND4_X1 _1994_ (
  .A1(_0254_),
  .A2(_0091_),
  .A3(_0098_),
  .A4(_0099_),
  .ZN(_0261_)
);

NAND3_X1 _1995_ (
  .A1(_0255_),
  .A2(_0260_),
  .A3(_0261_),
  .ZN(_0262_)
);

NAND2_X1 _1996_ (
  .A1(_0262_),
  .A2(_1125_),
  .ZN(_0263_)
);

INV_X1 _1997_ (
  .A(_1125_),
  .ZN(_0264_)
);

NAND4_X1 _1998_ (
  .A1(_0255_),
  .A2(_0260_),
  .A3(_0264_),
  .A4(_0261_),
  .ZN(_0265_)
);

NAND3_X1 _1999_ (
  .A1(_0263_),
  .A2(_0265_),
  .A3(_0584_),
  .ZN(_0266_)
);

NAND2_X1 _2000_ (
  .A1(_0581_),
  .A2(\ext_mult_res[18] ),
  .ZN(_0267_)
);

NAND2_X1 _2001_ (
  .A1(_0267_),
  .A2(_0371_),
  .ZN(_0268_)
);

INV_X1 _2002_ (
  .A(_0268_),
  .ZN(_0269_)
);

AOI21_X1 _2003_ (
  .A(_0250_),
  .B1(_0266_),
  .B2(_0269_),
  .ZN(_0037_)
);

NOR2_X1 _2004_ (
  .A1(_0368_),
  .A2(result[19]),
  .ZN(_0270_)
);

NAND2_X1 _2005_ (
  .A1(_1123_),
  .A2(_1125_),
  .ZN(_0271_)
);

NOR2_X1 _2006_ (
  .A1(_0229_),
  .A2(_0271_),
  .ZN(_0272_)
);

AND2_X1 _2007_ (
  .A1(_0189_),
  .A2(_0272_),
  .ZN(_0273_)
);

NAND2_X1 _2008_ (
  .A1(_0115_),
  .A2(_0273_),
  .ZN(_0274_)
);

INV_X1 _2009_ (
  .A(_1124_),
  .ZN(_0275_)
);

OAI21_X1 _2010_ (
  .A(_0275_),
  .B1(_0264_),
  .B2(_0256_),
  .ZN(_0276_)
);

INV_X1 _2011_ (
  .A(_0276_),
  .ZN(_0277_)
);

OAI21_X1 _2012_ (
  .A(_0277_),
  .B1(_0238_),
  .B2(_0271_),
  .ZN(_0278_)
);

AOI21_X1 _2013_ (
  .A(_0278_),
  .B1(_0272_),
  .B2(_0194_),
  .ZN(_0279_)
);

NAND3_X1 _2014_ (
  .A1(_0118_),
  .A2(_0119_),
  .A3(_0273_),
  .ZN(_0280_)
);

NAND3_X1 _2015_ (
  .A1(_0274_),
  .A2(_0279_),
  .A3(_0280_),
  .ZN(_0281_)
);

NAND2_X1 _2016_ (
  .A1(_0281_),
  .A2(_1127_),
  .ZN(_0282_)
);

INV_X1 _2017_ (
  .A(_1127_),
  .ZN(_0283_)
);

NAND4_X1 _2018_ (
  .A1(_0274_),
  .A2(_0279_),
  .A3(_0283_),
  .A4(_0280_),
  .ZN(_0284_)
);

NAND3_X1 _2019_ (
  .A1(_0282_),
  .A2(_0284_),
  .A3(_0584_),
  .ZN(_0285_)
);

AOI21_X1 _2020_ (
  .A(_0270_),
  .B1(_0285_),
  .B2(_0269_),
  .ZN(_0038_)
);

NOR2_X1 _2021_ (
  .A1(_0368_),
  .A2(result[20]),
  .ZN(_0286_)
);

NAND2_X1 _2022_ (
  .A1(_1125_),
  .A2(_1127_),
  .ZN(_0287_)
);

NOR2_X1 _2023_ (
  .A1(_0252_),
  .A2(_0287_),
  .ZN(_0288_)
);

AND2_X1 _2024_ (
  .A1(_0208_),
  .A2(_0288_),
  .ZN(_0289_)
);

NAND2_X1 _2025_ (
  .A1(_0137_),
  .A2(_0289_),
  .ZN(_0290_)
);

INV_X1 _2026_ (
  .A(_1126_),
  .ZN(_0291_)
);

OAI21_X1 _2027_ (
  .A(_0291_),
  .B1(_0283_),
  .B2(_0275_),
  .ZN(_0292_)
);

INV_X1 _2028_ (
  .A(_0292_),
  .ZN(_0293_)
);

OAI21_X1 _2029_ (
  .A(_0293_),
  .B1(_0258_),
  .B2(_0287_),
  .ZN(_0294_)
);

AOI21_X1 _2030_ (
  .A(_0294_),
  .B1(_0288_),
  .B2(_0214_),
  .ZN(_0295_)
);

NAND3_X1 _2031_ (
  .A1(_0612_),
  .A2(_0140_),
  .A3(_0289_),
  .ZN(_0296_)
);

NAND3_X1 _2032_ (
  .A1(_0290_),
  .A2(_0295_),
  .A3(_0296_),
  .ZN(_0297_)
);

NAND2_X1 _2033_ (
  .A1(_0297_),
  .A2(_1129_),
  .ZN(_0298_)
);

INV_X1 _2034_ (
  .A(_1129_),
  .ZN(_0299_)
);

NAND4_X1 _2035_ (
  .A1(_0290_),
  .A2(_0295_),
  .A3(_0299_),
  .A4(_0296_),
  .ZN(_0300_)
);

NAND3_X1 _2036_ (
  .A1(_0298_),
  .A2(_0300_),
  .A3(_0584_),
  .ZN(_0301_)
);

AOI21_X1 _2037_ (
  .A(_0286_),
  .B1(_0301_),
  .B2(_0269_),
  .ZN(_0039_)
);

NAND2_X1 _2038_ (
  .A1(_1127_),
  .A2(_1129_),
  .ZN(_0302_)
);

NOR2_X1 _2039_ (
  .A1(_0271_),
  .A2(_0302_),
  .ZN(_0303_)
);

NAND2_X1 _2040_ (
  .A1(_0230_),
  .A2(_0303_),
  .ZN(_0304_)
);

INV_X1 _2041_ (
  .A(_0304_),
  .ZN(_0305_)
);

NAND2_X1 _2042_ (
  .A1(_0161_),
  .A2(_0305_),
  .ZN(_0306_)
);

INV_X1 _2043_ (
  .A(_0303_),
  .ZN(_0307_)
);

AOI21_X1 _2044_ (
  .A(_0307_),
  .B1(_0234_),
  .B2(_0238_),
  .ZN(_0308_)
);

INV_X1 _2045_ (
  .A(_1128_),
  .ZN(_0309_)
);

OAI21_X1 _2046_ (
  .A(_0309_),
  .B1(_0299_),
  .B2(_0291_),
  .ZN(_0310_)
);

INV_X1 _2047_ (
  .A(_0310_),
  .ZN(_0311_)
);

OAI21_X1 _2048_ (
  .A(_0311_),
  .B1(_0277_),
  .B2(_0302_),
  .ZN(_0312_)
);

NOR2_X1 _2049_ (
  .A1(_0308_),
  .A2(_0312_),
  .ZN(_0313_)
);

NOR2_X1 _2050_ (
  .A1(_0165_),
  .A2(_0304_),
  .ZN(_0314_)
);

NAND2_X1 _2051_ (
  .A1(_0623_),
  .A2(_0314_),
  .ZN(_0315_)
);

XOR2_X1 _2052_ (
  .A(\ext_mult_res[18] ),
  .B(result[21]),
  .Z(_0316_)
);

NAND4_X1 _2053_ (
  .A1(_0306_),
  .A2(_0313_),
  .A3(_0315_),
  .A4(_0316_),
  .ZN(_0317_)
);

NAND3_X1 _2054_ (
  .A1(_0306_),
  .A2(_0313_),
  .A3(_0315_),
  .ZN(_0318_)
);

INV_X1 _2055_ (
  .A(_0316_),
  .ZN(_0319_)
);

NAND2_X1 _2056_ (
  .A1(_0318_),
  .A2(_0319_),
  .ZN(_0320_)
);

NAND2_X1 _2057_ (
  .A1(_0317_),
  .A2(_0320_),
  .ZN(_0321_)
);

NAND2_X1 _2058_ (
  .A1(_0321_),
  .A2(_0594_),
  .ZN(_0322_)
);

NAND2_X1 _2059_ (
  .A1(_0322_),
  .A2(_0267_),
  .ZN(_0323_)
);

NAND2_X1 _2060_ (
  .A1(_0323_),
  .A2(_0372_),
  .ZN(_0324_)
);

NAND2_X1 _2061_ (
  .A1(_0387_),
  .A2(result[21]),
  .ZN(_0325_)
);

NAND2_X1 _2062_ (
  .A1(_0324_),
  .A2(_0325_),
  .ZN(_0040_)
);

FA_X1 _2063_ (
  .A(_0676_),
  .B(_0677_),
  .CI(_0678_),
  .CO(_0679_),
  .S(_0680_)
);

FA_X1 _2064_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0684_),
  .S(_0685_)
);

FA_X1 _2065_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0689_),
  .S(_0690_)
);

FA_X1 _2066_ (
  .A(_0690_),
  .B(_0684_),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0692_),
  .S(_0693_)
);

FA_X1 _2067_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0697_),
  .S(_0698_)
);

FA_X1 _2068_ (
  .A(_0698_),
  .B(_0699_),
  .CI(_0700_),
  .CO(_0701_),
  .S(_0702_)
);

FA_X1 _2069_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0706_),
  .S(_0707_)
);

FA_X1 _2070_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0711_),
  .S(_0712_)
);

FA_X1 _2071_ (
  .A(_0707_),
  .B(_0697_),
  .CI(_0712_),
  .CO(_0713_),
  .S(_0714_)
);

FA_X1 _2072_ (
  .A(_0715_),
  .B(_0716_),
  .CI(_0717_),
  .CO(_0718_),
  .S(_0719_)
);

FA_X1 _2073_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0723_),
  .S(_0724_)
);

FA_X1 _2074_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0728_),
  .S(_0729_)
);

FA_X1 _2075_ (
  .A(_0724_),
  .B(_0706_),
  .CI(_0729_),
  .CO(_0730_),
  .S(_0731_)
);

FA_X1 _2076_ (
  .A(_0731_),
  .B(_0713_),
  .CI(_0732_),
  .CO(_0733_),
  .S(_0734_)
);

FA_X1 _2077_ (
  .A(_0735_),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0738_),
  .S(_0739_)
);

FA_X1 _2078_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0743_),
  .S(_0744_)
);

FA_X1 _2079_ (
  .A(_0744_),
  .B(_0739_),
  .CI(_0745_),
  .CO(_0746_),
  .S(_0747_)
);

FA_X1 _2080_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0751_),
  .S(_0752_)
);

FA_X1 _2081_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0756_),
  .S(_0757_)
);

FA_X1 _2082_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0761_),
  .S(_0762_)
);

FA_X1 _2083_ (
  .A(_0765_),
  .B(_0766_),
  .CI(_0767_),
  .CO(_0768_),
  .S(_0769_)
);

FA_X1 _2084_ (
  .A(_0770_),
  .B(_0747_),
  .CI(_0771_),
  .CO(_0772_),
  .S(_0773_)
);

FA_X1 _2085_ (
  .A(_0757_),
  .B(_0774_),
  .CI(_0775_),
  .CO(_0776_),
  .S(_0777_)
);

FA_X1 _2086_ (
  .A(_0778_),
  .B(_0779_),
  .CI(_0780_),
  .CO(_0781_),
  .S(_0782_)
);

FA_X1 _2087_ (
  .A(_0777_),
  .B(_0730_),
  .CI(_0784_),
  .CO(_0783_),
  .S(_0785_)
);

FA_X1 _2088_ (
  .A(_0786_),
  .B(_0733_),
  .CI(_0787_),
  .CO(_0788_),
  .S(_0789_)
);

FA_X1 _2089_ (
  .A(_0790_),
  .B(_0791_),
  .CI(_0792_),
  .CO(_0793_),
  .S(_0794_)
);

FA_X1 _2090_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(_0796_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0798_),
  .S(_0799_)
);

FA_X1 _2091_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0803_),
  .S(_0804_)
);

FA_X1 _2092_ (
  .A(_0799_),
  .B(_0738_),
  .CI(_0804_),
  .CO(_0805_),
  .S(_0806_)
);

FA_X1 _2093_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0809_),
  .S(_0810_)
);

FA_X1 _2094_ (
  .A(_0811_),
  .B(_0812_),
  .CI(_0813_),
  .CO(_0814_),
  .S(_0815_)
);

FA_X1 _2095_ (
  .A(_0806_),
  .B(_0746_),
  .CI(_0815_),
  .CO(_0816_),
  .S(_0817_)
);

FA_X1 _2096_ (
  .A(_0817_),
  .B(_0772_),
  .CI(_0818_),
  .CO(_0819_),
  .S(_0820_)
);

FA_X1 _2097_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(_0823_),
  .CO(_0824_),
  .S(_0825_)
);

FA_X1 _2098_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0829_),
  .S(_0830_)
);

FA_X1 _2099_ (
  .A(_0825_),
  .B(_0798_),
  .CI(_0830_),
  .CO(_0831_),
  .S(_0832_)
);

FA_X1 _2100_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0835_),
  .S(_0836_)
);

FA_X1 _2101_ (
  .A(_0837_),
  .B(_0838_),
  .CI(_0839_),
  .CO(_0840_),
  .S(_0841_)
);

FA_X1 _2102_ (
  .A(_0841_),
  .B(_0832_),
  .CI(_0805_),
  .CO(_0842_),
  .S(_0843_)
);

FA_X1 _2103_ (
  .A(_0816_),
  .B(_0843_),
  .CI(_0844_),
  .CO(_0845_),
  .S(_0846_)
);

FA_X1 _2104_ (
  .A(_0847_),
  .B(_0848_),
  .CI(_0849_),
  .CO(_0850_),
  .S(_0851_)
);

FA_X1 _2105_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0855_),
  .S(_0856_)
);

FA_X1 _2106_ (
  .A(_0857_),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0860_),
  .S(_0861_)
);

FA_X1 _2107_ (
  .A(_0862_),
  .B(_0824_),
  .CI(_0861_),
  .CO(_0863_),
  .S(_0864_)
);

FA_X1 _2108_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0867_),
  .S(_0868_)
);

FA_X1 _2109_ (
  .A(_0829_),
  .B(_0868_),
  .CI(_0835_),
  .CO(_0869_),
  .S(_0870_)
);

FA_X1 _2110_ (
  .A(_0864_),
  .B(_0831_),
  .CI(_0870_),
  .CO(_0871_),
  .S(_0872_)
);

FA_X1 _2111_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0874_),
  .S(_0875_)
);

FA_X1 _2112_ (
  .A(_0872_),
  .B(_0842_),
  .CI(_0876_),
  .CO(_0877_),
  .S(_0878_)
);

FA_X1 _2113_ (
  .A(_0878_),
  .B(_0845_),
  .CI(_0879_),
  .CO(_0880_),
  .S(_0881_)
);

FA_X1 _2114_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0883_),
  .S(_0884_)
);

FA_X1 _2115_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(_0886_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0888_),
  .S(_0889_)
);

FA_X1 _2116_ (
  .A(_0890_),
  .B(_0891_),
  .CI(_0889_),
  .CO(_0892_),
  .S(_0893_)
);

FA_X1 _2117_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0896_),
  .S(_0897_)
);

FA_X1 _2118_ (
  .A(_0860_),
  .B(_0897_),
  .CI(_0867_),
  .CO(_0898_),
  .S(_0899_)
);

FA_X1 _2119_ (
  .A(_0893_),
  .B(_0863_),
  .CI(_0899_),
  .CO(_0900_),
  .S(_0901_)
);

FA_X1 _2120_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0902_),
  .S(_0903_)
);

FA_X1 _2121_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(_0904_),
  .CI(_0905_),
  .CO(_0906_),
  .S(_0907_)
);

FA_X1 _2122_ (
  .A(_0908_),
  .B(_0909_),
  .CI(_0910_),
  .CO(_0911_),
  .S(_0912_)
);

FA_X1 _2123_ (
  .A(_0901_),
  .B(_0871_),
  .CI(_0913_),
  .CO(_0914_),
  .S(_0915_)
);

FA_X1 _2124_ (
  .A(_0915_),
  .B(_0877_),
  .CI(_0916_),
  .CO(_0917_),
  .S(_0918_)
);

FA_X1 _2125_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(_0921_),
  .CO(_0922_),
  .S(_0923_)
);

FA_X1 _2126_ (
  .A(_0924_),
  .B(_0923_),
  .CI(_0890_),
  .CO(_0925_),
  .S(_0926_)
);

FA_X1 _2127_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0929_),
  .S(_0930_)
);

FA_X1 _2128_ (
  .A(_0888_),
  .B(_0930_),
  .CI(_0896_),
  .CO(_0931_),
  .S(_0932_)
);

FA_X1 _2129_ (
  .A(_0926_),
  .B(_0892_),
  .CI(_0932_),
  .CO(_0933_),
  .S(_0934_)
);

FA_X1 _2130_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0935_),
  .S(_0936_)
);

FA_X1 _2131_ (
  .A(_0937_),
  .B(_0938_),
  .CI(_0902_),
  .CO(_0939_),
  .S(_0940_)
);

FA_X1 _2132_ (
  .A(_0898_),
  .B(_0940_),
  .CI(_0906_),
  .CO(_0943_),
  .S(_0944_)
);

FA_X1 _2133_ (
  .A(_0934_),
  .B(_0900_),
  .CI(_0944_),
  .CO(_0945_),
  .S(_0946_)
);

FA_X1 _2134_ (
  .A(_0947_),
  .B(_0948_),
  .CI(_0911_),
  .CO(_0949_),
  .S(_0950_)
);

FA_X1 _2135_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0954_),
  .S(_0955_)
);

FA_X1 _2136_ (
  .A(_0924_),
  .B(_0956_),
  .CI(_0890_),
  .CO(_0957_),
  .S(_0958_)
);

FA_X1 _2137_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(_0959_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0961_),
  .S(_0962_)
);

FA_X1 _2138_ (
  .A(_0922_),
  .B(_0962_),
  .CI(_0929_),
  .CO(_0963_),
  .S(_0964_)
);

FA_X1 _2139_ (
  .A(_0958_),
  .B(_0925_),
  .CI(_0964_),
  .CO(_0965_),
  .S(_0966_)
);

FA_X1 _2140_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0967_),
  .S(_0968_)
);

FA_X1 _2141_ (
  .A(_0969_),
  .B(_0970_),
  .CI(_0935_),
  .CO(_0971_),
  .S(_0972_)
);

FA_X1 _2142_ (
  .A(_0974_),
  .B(_0975_),
  .CI(_0976_),
  .CO(_0977_),
  .S(_0978_)
);

FA_X1 _2143_ (
  .A(_0966_),
  .B(_0933_),
  .CI(_0978_),
  .CO(_0979_),
  .S(_0980_)
);

FA_X1 _2144_ (
  .A(_0981_),
  .B(_0982_),
  .CI(_0983_),
  .CO(_0984_),
  .S(_0985_)
);

FA_X1 _2145_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0987_),
  .S(_0988_)
);

FA_X1 _2146_ (
  .A(_0924_),
  .B(_0989_),
  .CI(_0890_),
  .CO(_0990_),
  .S(_0991_)
);

FA_X1 _2147_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(_0993_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0994_),
  .S(_0995_)
);

FA_X1 _2148_ (
  .A(_0995_),
  .B(_0961_),
  .CI(_0996_),
  .CO(_0997_),
  .S(_0998_)
);

FA_X1 _2149_ (
  .A(_0998_),
  .B(_0991_),
  .CI(_0957_),
  .CO(_0999_),
  .S(_1000_)
);

FA_X1 _2150_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_1004_),
  .S(_1005_)
);

FA_X1 _2151_ (
  .A(_1005_),
  .B(_1006_),
  .CI(_0903_),
  .CO(_1007_),
  .S(_1008_)
);

FA_X1 _2152_ (
  .A(_1009_),
  .B(_1008_),
  .CI(_1010_),
  .CO(_1011_),
  .S(_1012_)
);

FA_X1 _2153_ (
  .A(_1000_),
  .B(_0965_),
  .CI(_1012_),
  .CO(_1013_),
  .S(_1014_)
);

FA_X1 _2154_ (
  .A(_1014_),
  .B(_0979_),
  .CI(_1015_),
  .CO(_1016_),
  .S(_1017_)
);

FA_X1 _2155_ (
  .A(_1018_),
  .B(_0984_),
  .CI(_1019_),
  .CO(_1020_),
  .S(_1021_)
);

FA_X1 _2156_ (
  .A(_1022_),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_1025_),
  .S(_1026_)
);

FA_X1 _2157_ (
  .A(_1027_),
  .B(_1028_),
  .CI(_0994_),
  .CO(_1029_),
  .S(_1030_)
);

FA_X1 _2158_ (
  .A(_0990_),
  .B(_1030_),
  .CI(_0991_),
  .CO(_1031_),
  .S(_1032_)
);

FA_X1 _2159_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_1034_),
  .S(_1035_)
);

FA_X1 _2160_ (
  .A(_1035_),
  .B(_1004_),
  .CI(_0936_),
  .CO(_1036_),
  .S(_1037_)
);

FA_X1 _2161_ (
  .A(_0997_),
  .B(_1038_),
  .CI(_1039_),
  .CO(_1040_),
  .S(_1041_)
);

FA_X1 _2162_ (
  .A(_1032_),
  .B(_0999_),
  .CI(_1041_),
  .CO(_1042_),
  .S(_1043_)
);

FA_X1 _2163_ (
  .A(_1043_),
  .B(_1013_),
  .CI(_1044_),
  .CO(_1045_),
  .S(_1046_)
);

FA_X1 _2164_ (
  .A(_1047_),
  .B(_1048_),
  .CI(_1049_),
  .CO(_1050_),
  .S(_1051_)
);

FA_X1 _2165_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_1055_),
  .S(_1056_)
);

FA_X1 _2166_ (
  .A(_1027_),
  .B(_1057_),
  .CI(_1058_),
  .CO(_1059_),
  .S(_1060_)
);

FA_X1 _2167_ (
  .A(_0990_),
  .B(_1060_),
  .CI(_0991_),
  .CO(_1061_),
  .S(_1062_)
);

FA_X1 _2168_ (
  .A(_0993_),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_1063_),
  .S(_1064_)
);

FA_X1 _2169_ (
  .A(_1034_),
  .B(_1064_),
  .CI(_0968_),
  .CO(_1065_),
  .S(_1066_)
);

FA_X1 _2170_ (
  .A(_1066_),
  .B(_1036_),
  .CI(_1067_),
  .CO(_1068_),
  .S(_1069_)
);

FA_X1 _2171_ (
  .A(_1069_),
  .B(_1062_),
  .CI(_1031_),
  .CO(_1070_),
  .S(_1071_)
);

FA_X1 _2172_ (
  .A(_0973_),
  .B(_0875_),
  .CI(_1072_),
  .CO(_1073_),
  .S(_1074_)
);

FA_X1 _2173_ (
  .A(_1075_),
  .B(_1076_),
  .CI(_1077_),
  .CO(_1078_),
  .S(_1079_)
);

FA_X1 _2174_ (
  .A(_1071_),
  .B(_1042_),
  .CI(_1080_),
  .CO(_1081_),
  .S(_1082_)
);

FA_X1 _2175_ (
  .A(_1083_),
  .B(_1084_),
  .CI(_1085_),
  .CO(_1086_),
  .S(_1087_)
);

HA_X1 _2176_ (
  .A(result[0]),
  .B(\ext_mult_res[0] ),
  .CO(_1088_),
  .S(_1089_)
);

HA_X1 _2177_ (
  .A(result[1]),
  .B(\ext_mult_res[1] ),
  .CO(_1090_),
  .S(_1091_)
);

HA_X1 _2178_ (
  .A(result[2]),
  .B(\ext_mult_res[2] ),
  .CO(_1092_),
  .S(_1093_)
);

HA_X1 _2179_ (
  .A(result[3]),
  .B(\ext_mult_res[3] ),
  .CO(_1094_),
  .S(_1095_)
);

HA_X1 _2180_ (
  .A(result[4]),
  .B(\ext_mult_res[4] ),
  .CO(_1096_),
  .S(_1097_)
);

HA_X1 _2181_ (
  .A(result[5]),
  .B(\ext_mult_res[5] ),
  .CO(_1098_),
  .S(_1099_)
);

HA_X1 _2182_ (
  .A(result[6]),
  .B(\ext_mult_res[6] ),
  .CO(_1100_),
  .S(_1101_)
);

HA_X1 _2183_ (
  .A(result[7]),
  .B(\ext_mult_res[7] ),
  .CO(_1102_),
  .S(_1103_)
);

HA_X1 _2184_ (
  .A(result[8]),
  .B(\ext_mult_res[8] ),
  .CO(_1104_),
  .S(_1105_)
);

HA_X1 _2185_ (
  .A(result[9]),
  .B(\ext_mult_res[9] ),
  .CO(_1106_),
  .S(_1107_)
);

HA_X1 _2186_ (
  .A(result[10]),
  .B(\ext_mult_res[10] ),
  .CO(_1108_),
  .S(_1109_)
);

HA_X1 _2187_ (
  .A(result[11]),
  .B(\ext_mult_res[11] ),
  .CO(_1110_),
  .S(_1111_)
);

HA_X1 _2188_ (
  .A(result[12]),
  .B(\ext_mult_res[12] ),
  .CO(_1112_),
  .S(_1113_)
);

HA_X1 _2189_ (
  .A(result[13]),
  .B(\ext_mult_res[13] ),
  .CO(_1114_),
  .S(_1115_)
);

HA_X1 _2190_ (
  .A(result[14]),
  .B(\ext_mult_res[14] ),
  .CO(_1116_),
  .S(_1117_)
);

HA_X1 _2191_ (
  .A(result[15]),
  .B(\ext_mult_res[15] ),
  .CO(_1118_),
  .S(_1119_)
);

HA_X1 _2192_ (
  .A(result[16]),
  .B(\ext_mult_res[16] ),
  .CO(_1120_),
  .S(_1121_)
);

HA_X1 _2193_ (
  .A(result[17]),
  .B(\ext_mult_res[17] ),
  .CO(_1122_),
  .S(_1123_)
);

HA_X1 _2194_ (
  .A(result[18]),
  .B(\ext_mult_res[18] ),
  .CO(_1124_),
  .S(_1125_)
);

HA_X1 _2195_ (
  .A(result[19]),
  .B(\ext_mult_res[18] ),
  .CO(_1126_),
  .S(_1127_)
);

HA_X1 _2196_ (
  .A(result[20]),
  .B(\ext_mult_res[18] ),
  .CO(_1128_),
  .S(_1129_)
);

HA_X1 _2197_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_1132_),
  .S(_1133_)
);

HA_X1 _2198_ (
  .A(_0685_),
  .B(_1132_),
  .CO(_1134_),
  .S(_1135_)
);

HA_X1 _2199_ (
  .A(_0693_),
  .B(_1134_),
  .CO(_1136_),
  .S(_1137_)
);

HA_X1 _2200_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0717_),
  .S(_1140_)
);

HA_X1 _2201_ (
  .A(_1141_),
  .B(_0692_),
  .CO(_1142_),
  .S(_1143_)
);

HA_X1 _2202_ (
  .A(_1143_),
  .B(_1136_),
  .CO(_1144_),
  .S(_1145_)
);

HA_X1 _2203_ (
  .A(_0719_),
  .B(_1142_),
  .CO(_1146_),
  .S(_1147_)
);

HA_X1 _2204_ (
  .A(_1147_),
  .B(_1144_),
  .CO(_1148_),
  .S(_1149_)
);

HA_X1 _2205_ (
  .A(_1150_),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_1152_),
  .S(_1153_)
);

HA_X1 _2206_ (
  .A(_1154_),
  .B(_0718_),
  .CO(_1155_),
  .S(_1156_)
);

HA_X1 _2207_ (
  .A(_1156_),
  .B(_1146_),
  .CO(_1157_),
  .S(_1158_)
);

HA_X1 _2208_ (
  .A(_1158_),
  .B(_1148_),
  .CO(_1159_),
  .S(_1160_)
);

HA_X1 _2209_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_0767_),
  .S(_1162_)
);

HA_X1 _2210_ (
  .A(_1163_),
  .B(_1162_),
  .CO(_0780_),
  .S(_1164_)
);

HA_X1 _2211_ (
  .A(_0782_),
  .B(_1165_),
  .CO(_1166_),
  .S(_1167_)
);

HA_X1 _2212_ (
  .A(_1167_),
  .B(_1168_),
  .CO(_1169_),
  .S(_1170_)
);

HA_X1 _2213_ (
  .A(_1171_),
  .B(_1155_),
  .CO(_1168_),
  .S(_1172_)
);

HA_X1 _2214_ (
  .A(_1170_),
  .B(_1173_),
  .CO(_1174_),
  .S(_1175_)
);

HA_X1 _2215_ (
  .A(_1172_),
  .B(_1157_),
  .CO(_1173_),
  .S(_1176_)
);

HA_X1 _2216_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(_0768_),
  .CO(_0847_),
  .S(_1178_)
);

HA_X1 _2217_ (
  .A(_1179_),
  .B(_0781_),
  .CO(_1180_),
  .S(_1181_)
);

HA_X1 _2218_ (
  .A(_1181_),
  .B(_1166_),
  .CO(_1182_),
  .S(_1183_)
);

HA_X1 _2219_ (
  .A(_1183_),
  .B(_1169_),
  .CO(_1184_),
  .S(_1185_)
);

HA_X1 _2220_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .CO(_1072_),
  .S(_0941_)
);

HA_X1 _2221_ (
  .A(_0814_),
  .B(_0941_),
  .CO(_1186_),
  .S(_1187_)
);

HA_X1 _2222_ (
  .A(_0851_),
  .B(_1180_),
  .CO(_1188_),
  .S(_1189_)
);

HA_X1 _2223_ (
  .A(_1189_),
  .B(_1182_),
  .CO(_1190_),
  .S(_1191_)
);

HA_X1 _2224_ (
  .A(_0875_),
  .B(_1072_),
  .CO(_0910_),
  .S(_1192_)
);

HA_X1 _2225_ (
  .A(_0840_),
  .B(_1192_),
  .CO(_1193_),
  .S(_1194_)
);

HA_X1 _2226_ (
  .A(_0881_),
  .B(_0850_),
  .CO(_1195_),
  .S(_1196_)
);

HA_X1 _2227_ (
  .A(_1196_),
  .B(_1188_),
  .CO(_1197_),
  .S(_1198_)
);

HA_X1 _2228_ (
  .A(_1199_),
  .B(_0918_),
  .CO(_1200_),
  .S(_1201_)
);

HA_X1 _2229_ (
  .A(_1195_),
  .B(_1201_),
  .CO(_1202_),
  .S(_1203_)
);

HA_X1 _2230_ (
  .A(_1204_),
  .B(_1205_),
  .CO(_1206_),
  .S(_1207_)
);

HA_X1 _2231_ (
  .A(_1207_),
  .B(_1200_),
  .CO(_1208_),
  .S(_1209_)
);

HA_X1 _2232_ (
  .A(_1210_),
  .B(_1072_),
  .CO(_1019_),
  .S(_0981_)
);

HA_X1 _2233_ (
  .A(_1211_),
  .B(_0949_),
  .CO(_1212_),
  .S(_1213_)
);

HA_X1 _2234_ (
  .A(_1213_),
  .B(_1206_),
  .CO(_1214_),
  .S(_1215_)
);

HA_X1 _2235_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 ),
  .B(_0874_),
  .CO(_1217_),
  .S(_1218_)
);

HA_X1 _2236_ (
  .A(_0977_),
  .B(_1218_),
  .CO(_1049_),
  .S(_1219_)
);

HA_X1 _2237_ (
  .A(_1021_),
  .B(_1212_),
  .CO(_1220_),
  .S(_1221_)
);

HA_X1 _2238_ (
  .A(_1222_),
  .B(_1216_),
  .CO(_1223_),
  .S(_1224_)
);

HA_X1 _2239_ (
  .A(_0941_),
  .B(_0942_),
  .CO(_1225_),
  .S(_1226_)
);

HA_X1 _2240_ (
  .A(_1226_),
  .B(_1217_),
  .CO(_1077_),
  .S(_1227_)
);

HA_X1 _2241_ (
  .A(_1011_),
  .B(_1227_),
  .CO(_1085_),
  .S(_1228_)
);

HA_X1 _2242_ (
  .A(_1051_),
  .B(_1020_),
  .CO(_1229_),
  .S(_1230_)
);

HA_X1 _2243_ (
  .A(_1074_),
  .B(_1225_),
  .CO(_1231_),
  .S(_1076_)
);

HA_X1 _2244_ (
  .A(_1087_),
  .B(_1050_),
  .CO(_1232_),
  .S(_1233_)
);

HA_X1 _2245_ (
  .A(_1176_),
  .B(_1159_),
  .CO(_1177_),
  .S(_1234_)
);

DFF_X1 \ext_mult_res[0]$_DFFE_PP_  (
  .D(_0000_),
  .CK(clk),
  .Q(\ext_mult_res[0] ),
  .QN(_0675_)
);

DFF_X1 \ext_mult_res[10]$_DFFE_PP_  (
  .D(_0010_),
  .CK(clk),
  .Q(\ext_mult_res[10] ),
  .QN(_0666_)
);

DFF_X1 \ext_mult_res[11]$_DFFE_PP_  (
  .D(_0011_),
  .CK(clk),
  .Q(\ext_mult_res[11] ),
  .QN(_0665_)
);

DFF_X1 \ext_mult_res[12]$_DFFE_PP_  (
  .D(_0012_),
  .CK(clk),
  .Q(\ext_mult_res[12] ),
  .QN(_0664_)
);

DFF_X1 \ext_mult_res[13]$_DFFE_PP_  (
  .D(_0013_),
  .CK(clk),
  .Q(\ext_mult_res[13] ),
  .QN(_0663_)
);

DFF_X1 \ext_mult_res[14]$_DFFE_PP_  (
  .D(_0014_),
  .CK(clk),
  .Q(\ext_mult_res[14] ),
  .QN(_0662_)
);

DFF_X1 \ext_mult_res[15]$_DFFE_PP_  (
  .D(_0015_),
  .CK(clk),
  .Q(\ext_mult_res[15] ),
  .QN(_0661_)
);

DFF_X1 \ext_mult_res[16]$_DFFE_PP_  (
  .D(_0016_),
  .CK(clk),
  .Q(\ext_mult_res[16] ),
  .QN(_0660_)
);

DFF_X1 \ext_mult_res[17]$_DFFE_PP_  (
  .D(_0017_),
  .CK(clk),
  .Q(\ext_mult_res[17] ),
  .QN(_0659_)
);

DFF_X1 \ext_mult_res[1]$_DFFE_PP_  (
  .D(_0001_),
  .CK(clk),
  .Q(\ext_mult_res[1] ),
  .QN(_0677_)
);

DFF_X1 \ext_mult_res[21]$_DFFE_PP_  (
  .D(_0018_),
  .CK(clk),
  .Q(\ext_mult_res[18] ),
  .QN(_0658_)
);

DFF_X1 \ext_mult_res[2]$_DFFE_PP_  (
  .D(_0002_),
  .CK(clk),
  .Q(\ext_mult_res[2] ),
  .QN(_0674_)
);

DFF_X1 \ext_mult_res[3]$_DFFE_PP_  (
  .D(_0003_),
  .CK(clk),
  .Q(\ext_mult_res[3] ),
  .QN(_0673_)
);

DFF_X1 \ext_mult_res[4]$_DFFE_PP_  (
  .D(_0004_),
  .CK(clk),
  .Q(\ext_mult_res[4] ),
  .QN(_0672_)
);

DFF_X1 \ext_mult_res[5]$_DFFE_PP_  (
  .D(_0005_),
  .CK(clk),
  .Q(\ext_mult_res[5] ),
  .QN(_0671_)
);

DFF_X1 \ext_mult_res[6]$_DFFE_PP_  (
  .D(_0006_),
  .CK(clk),
  .Q(\ext_mult_res[6] ),
  .QN(_0670_)
);

DFF_X1 \ext_mult_res[7]$_DFFE_PP_  (
  .D(_0007_),
  .CK(clk),
  .Q(\ext_mult_res[7] ),
  .QN(_0669_)
);

DFF_X1 \ext_mult_res[8]$_DFFE_PP_  (
  .D(_0008_),
  .CK(clk),
  .Q(\ext_mult_res[8] ),
  .QN(_0668_)
);

DFF_X1 \ext_mult_res[9]$_DFFE_PP_  (
  .D(_0009_),
  .CK(clk),
  .Q(\ext_mult_res[9] ),
  .QN(_0667_)
);

DFF_X1 \result[0]$_DFFE_PP_  (
  .D(_0019_),
  .CK(clk),
  .Q(result[0]),
  .QN(_0657_)
);

DFF_X1 \result[10]$_DFFE_PP_  (
  .D(_0029_),
  .CK(clk),
  .Q(result[10]),
  .QN(_0648_)
);

DFF_X1 \result[11]$_DFFE_PP_  (
  .D(_0030_),
  .CK(clk),
  .Q(result[11]),
  .QN(_0647_)
);

DFF_X1 \result[12]$_DFFE_PP_  (
  .D(_0031_),
  .CK(clk),
  .Q(result[12]),
  .QN(_0646_)
);

DFF_X1 \result[13]$_DFFE_PP_  (
  .D(_0032_),
  .CK(clk),
  .Q(result[13]),
  .QN(_0645_)
);

DFF_X1 \result[14]$_DFFE_PP_  (
  .D(_0033_),
  .CK(clk),
  .Q(result[14]),
  .QN(_0644_)
);

DFF_X1 \result[15]$_DFFE_PP_  (
  .D(_0034_),
  .CK(clk),
  .Q(result[15]),
  .QN(_0643_)
);

DFF_X1 \result[16]$_DFFE_PP_  (
  .D(_0035_),
  .CK(clk),
  .Q(result[16]),
  .QN(_0642_)
);

DFF_X1 \result[17]$_DFFE_PP_  (
  .D(_0036_),
  .CK(clk),
  .Q(result[17]),
  .QN(_0641_)
);

DFF_X1 \result[18]$_DFFE_PP_  (
  .D(_0037_),
  .CK(clk),
  .Q(result[18]),
  .QN(_0640_)
);

DFF_X1 \result[19]$_DFFE_PP_  (
  .D(_0038_),
  .CK(clk),
  .Q(result[19]),
  .QN(_0639_)
);

DFF_X1 \result[1]$_DFFE_PP_  (
  .D(_0020_),
  .CK(clk),
  .Q(result[1]),
  .QN(_0676_)
);

DFF_X1 \result[20]$_DFFE_PP_  (
  .D(_0039_),
  .CK(clk),
  .Q(result[20]),
  .QN(_0638_)
);

DFF_X1 \result[21]$_DFFE_PP_  (
  .D(_0040_),
  .CK(clk),
  .Q(result[21]),
  .QN(_0637_)
);

DFF_X1 \result[2]$_DFFE_PP_  (
  .D(_0021_),
  .CK(clk),
  .Q(result[2]),
  .QN(_0656_)
);

DFF_X1 \result[3]$_DFFE_PP_  (
  .D(_0022_),
  .CK(clk),
  .Q(result[3]),
  .QN(_0655_)
);

DFF_X1 \result[4]$_DFFE_PP_  (
  .D(_0023_),
  .CK(clk),
  .Q(result[4]),
  .QN(_0654_)
);

DFF_X1 \result[5]$_DFFE_PP_  (
  .D(_0024_),
  .CK(clk),
  .Q(result[5]),
  .QN(_0653_)
);

DFF_X1 \result[6]$_DFFE_PP_  (
  .D(_0025_),
  .CK(clk),
  .Q(result[6]),
  .QN(_0652_)
);

DFF_X1 \result[7]$_DFFE_PP_  (
  .D(_0026_),
  .CK(clk),
  .Q(result[7]),
  .QN(_0651_)
);

DFF_X1 \result[8]$_DFFE_PP_  (
  .D(_0027_),
  .CK(clk),
  .Q(result[8]),
  .QN(_0650_)
);

DFF_X1 \result[9]$_DFFE_PP_  (
  .D(_0028_),
  .CK(clk),
  .Q(result[9]),
  .QN(_0649_)
);

LOGIC0_X1 \logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002  (
  .Z(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 )
);

LOGIC1_X1 \logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002  (
  .Z(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002 )
);

INV_X1 _1283__reduced (
  .A(_0326_),
  .ZN(_0735_)
);

INV_X1 _1308__reduced (
  .A(_0333_),
  .ZN(_0796_)
);

INV_X1 _1319__reduced (
  .A(_0339_),
  .ZN(_0823_)
);

INV_X1 _1328__reduced (
  .A(_0341_),
  .ZN(_0857_)
);

INV_X1 _1337__reduced (
  .A(_0354_),
  .ZN(_0886_)
);

INV_X1 _1345__reduced (
  .A(_0355_),
  .ZN(_0921_)
);

INV_X1 _1353__reduced (
  .A(_0348_),
  .ZN(_0959_)
);

INV_X1 _1359__reduced (
  .A(din[7]),
  .ZN(_0993_)
);

NOR2_X1 _1473__reduced (
  .A1(_0370_),
  .A2(_0372_),
  .ZN(_0000_)
);

NAND2_X1 _1619__reduced (
  .A1(_0497_),
  .A2(_0498_),
  .ZN(_0501_)
);

INV_X1 _1620__reduced (
  .A(_0501_),
  .ZN(_0502_)
);

INV_X1 _1634__reduced (
  .A(_0993_),
  .ZN(_0516_)
);

INV_X1 _1636__reduced (
  .A(_0516_),
  .ZN(_0518_)
);

INV_X1 _1637__reduced (
  .A(_0518_),
  .ZN(_0519_)
);

INV_X1 _1639__reduced (
  .A(_0519_),
  .ZN(_0521_)
);

INV_X1 _1643__reduced (
  .A(_0516_),
  .ZN(_0525_)
);

INV_X1 _1644__reduced (
  .A(_0525_),
  .ZN(_0526_)
);

NAND2_X1 _1662__reduced (
  .A1(_0540_),
  .A2(_0541_),
  .ZN(_0544_)
);

INV_X1 _1663__reduced (
  .A(_0544_),
  .ZN(_0545_)
);

NAND2_X1 _1667__reduced (
  .A1(_0544_),
  .A2(_0546_),
  .ZN(_0549_)
);
endmodule //$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002

module \$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 (input clk,
 input ena, input dclr, input [7:0] din, input [10:0] coef, output [21:0] result);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire _0032_;
wire _0033_;
wire _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire _0066_;
wire _0067_;
wire _0068_;
wire _0069_;
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0333_;
wire _0339_;
wire _0341_;
wire _0348_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0367_;
wire _0368_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
wire _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
wire _0444_;
wire _0445_;
wire _0446_;
wire _0447_;
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire _0658_;
wire _0659_;
wire _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire _0673_;
wire _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire _0679_;
wire _0680_;
wire _0684_;
wire _0685_;
wire _0689_;
wire _0690_;
wire _0692_;
wire _0693_;
wire _0697_;
wire _0698_;
wire _0699_;
wire _0700_;
wire _0701_;
wire _0702_;
wire _0706_;
wire _0707_;
wire _0711_;
wire _0712_;
wire _0713_;
wire _0714_;
wire _0715_;
wire _0716_;
wire _0717_;
wire _0718_;
wire _0719_;
wire _0723_;
wire _0724_;
wire _0728_;
wire _0729_;
wire _0730_;
wire _0731_;
wire _0732_;
wire _0733_;
wire _0734_;
wire _0735_;
wire _0738_;
wire _0739_;
wire _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0751_;
wire _0752_;
wire _0756_;
wire _0757_;
wire _0761_;
wire _0762_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire _0780_;
wire _0781_;
wire _0782_;
wire _0783_;
wire _0784_;
wire _0785_;
wire _0786_;
wire _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire _0795_;
wire _0796_;
wire _0798_;
wire _0799_;
wire _0803_;
wire _0804_;
wire _0805_;
wire _0806_;
wire _0809_;
wire _0810_;
wire _0811_;
wire _0812_;
wire _0813_;
wire _0814_;
wire _0815_;
wire _0816_;
wire _0817_;
wire _0818_;
wire _0819_;
wire _0820_;
wire _0821_;
wire _0822_;
wire _0823_;
wire _0824_;
wire _0825_;
wire _0829_;
wire _0830_;
wire _0831_;
wire _0832_;
wire _0835_;
wire _0836_;
wire _0837_;
wire _0838_;
wire _0839_;
wire _0840_;
wire _0841_;
wire _0842_;
wire _0843_;
wire _0844_;
wire _0845_;
wire _0846_;
wire _0847_;
wire _0848_;
wire _0849_;
wire _0850_;
wire _0851_;
wire _0852_;
wire _0853_;
wire _0854_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0860_;
wire _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0867_;
wire _0868_;
wire _0869_;
wire _0870_;
wire _0871_;
wire _0872_;
wire _0874_;
wire _0875_;
wire _0876_;
wire _0877_;
wire _0878_;
wire _0879_;
wire _0880_;
wire _0881_;
wire _0882_;
wire _0883_;
wire _0884_;
wire _0885_;
wire _0886_;
wire _0888_;
wire _0889_;
wire _0890_;
wire _0891_;
wire _0892_;
wire _0893_;
wire _0896_;
wire _0897_;
wire _0898_;
wire _0899_;
wire _0900_;
wire _0901_;
wire _0902_;
wire _0903_;
wire _0904_;
wire _0905_;
wire _0906_;
wire _0907_;
wire _0908_;
wire _0909_;
wire _0910_;
wire _0911_;
wire _0912_;
wire _0913_;
wire _0914_;
wire _0915_;
wire _0916_;
wire _0917_;
wire _0918_;
wire _0919_;
wire _0920_;
wire _0921_;
wire _0922_;
wire _0923_;
wire _0924_;
wire _0925_;
wire _0926_;
wire _0929_;
wire _0930_;
wire _0931_;
wire _0932_;
wire _0933_;
wire _0934_;
wire _0935_;
wire _0936_;
wire _0937_;
wire _0938_;
wire _0939_;
wire _0940_;
wire _0941_;
wire _0942_;
wire _0943_;
wire _0944_;
wire _0945_;
wire _0946_;
wire _0947_;
wire _0948_;
wire _0949_;
wire _0950_;
wire _0951_;
wire _0952_;
wire _0953_;
wire _0954_;
wire _0955_;
wire _0956_;
wire _0957_;
wire _0958_;
wire _0959_;
wire _0961_;
wire _0962_;
wire _0963_;
wire _0964_;
wire _0965_;
wire _0966_;
wire _0967_;
wire _0968_;
wire _0969_;
wire _0970_;
wire _0971_;
wire _0972_;
wire _0973_;
wire _0974_;
wire _0975_;
wire _0976_;
wire _0977_;
wire _0978_;
wire _0979_;
wire _0980_;
wire _0981_;
wire _0982_;
wire _0983_;
wire _0984_;
wire _0985_;
wire _0986_;
wire _0987_;
wire _0988_;
wire _0989_;
wire _0990_;
wire _0991_;
wire _0992_;
wire _0993_;
wire _0994_;
wire _0995_;
wire _0996_;
wire _0997_;
wire _0998_;
wire _0999_;
wire _1000_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire \ext_mult_res[0] ;
wire \ext_mult_res[10] ;
wire \ext_mult_res[11] ;
wire \ext_mult_res[12] ;
wire \ext_mult_res[13] ;
wire \ext_mult_res[14] ;
wire \ext_mult_res[15] ;
wire \ext_mult_res[16] ;
wire \ext_mult_res[17] ;
wire \ext_mult_res[18] ;
wire \ext_mult_res[1] ;
wire \ext_mult_res[2] ;
wire \ext_mult_res[3] ;
wire \ext_mult_res[4] ;
wire \ext_mult_res[5] ;
wire \ext_mult_res[6] ;
wire \ext_mult_res[7] ;
wire \ext_mult_res[8] ;
wire \ext_mult_res[9] ;
wire \logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ;
wire \logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ;

BUF_X1 _1235_ (
  .A(din[0]),
  .Z(_0326_)
);

BUF_X1 _1245_ (
  .A(din[1]),
  .Z(_0333_)
);

BUF_X1 _1255_ (
  .A(din[2]),
  .Z(_0339_)
);

BUF_X1 _1258_ (
  .A(din[3]),
  .Z(_0341_)
);

BUF_X1 _1279_ (
  .A(din[6]),
  .Z(_0348_)
);

BUF_X1 _1292_ (
  .A(din[4]),
  .Z(_0354_)
);

BUF_X1 _1294_ (
  .A(din[5]),
  .Z(_0355_)
);

BUF_X8 _1299_ (
  .A(din[7]),
  .Z(_0356_)
);

BUF_X4 _1306_ (
  .A(coef[9]),
  .Z(_0358_)
);

NAND2_X1 _1307_ (
  .A1(_0326_),
  .A2(_0358_),
  .ZN(_0795_)
);

BUF_X4 _1316_ (
  .A(coef[10]),
  .Z(_0359_)
);

NAND2_X1 _1317_ (
  .A1(_0326_),
  .A2(_0359_),
  .ZN(_0821_)
);

INV_X1 _1318_ (
  .A(_0821_),
  .ZN(_0854_)
);

NAND2_X1 _1324_ (
  .A1(_0333_),
  .A2(_0359_),
  .ZN(_0360_)
);

INV_X1 _1325_ (
  .A(_0360_),
  .ZN(_0852_)
);

NAND2_X1 _1326_ (
  .A1(_0339_),
  .A2(_0358_),
  .ZN(_0361_)
);

INV_X1 _1327_ (
  .A(_0361_),
  .ZN(_0853_)
);

NAND2_X1 _1334_ (
  .A1(_0339_),
  .A2(_0359_),
  .ZN(_0362_)
);

INV_X1 _1335_ (
  .A(_0362_),
  .ZN(_0882_)
);

NAND2_X1 _1336_ (
  .A1(_0341_),
  .A2(_0358_),
  .ZN(_0885_)
);

INV_X1 _1342_ (
  .A(_1177_),
  .ZN(_0792_)
);

NAND2_X1 _1343_ (
  .A1(din[3]),
  .A2(_0359_),
  .ZN(_0919_)
);

INV_X1 _1344_ (
  .A(_0919_),
  .ZN(_0951_)
);

NAND2_X1 _1349_ (
  .A1(_0354_),
  .A2(_0359_),
  .ZN(_0363_)
);

INV_X1 _1350_ (
  .A(_0363_),
  .ZN(_0952_)
);

NAND2_X1 _1351_ (
  .A1(din[5]),
  .A2(_0358_),
  .ZN(_0364_)
);

INV_X1 _1352_ (
  .A(_0364_),
  .ZN(_0953_)
);

NAND2_X1 _1356_ (
  .A1(_0355_),
  .A2(_0359_),
  .ZN(_0365_)
);

INV_X1 _1357_ (
  .A(_0365_),
  .ZN(_0986_)
);

NAND2_X1 _1358_ (
  .A1(_0348_),
  .A2(_0358_),
  .ZN(_0992_)
);

INV_X1 _1360_ (
  .A(_0993_),
  .ZN(_1022_)
);

NAND2_X2 _1361_ (
  .A1(din[6]),
  .A2(_0359_),
  .ZN(_1052_)
);

INV_X2 _1362_ (
  .A(_1052_),
  .ZN(_1023_)
);

NAND2_X2 _1363_ (
  .A1(_0356_),
  .A2(_0358_),
  .ZN(_1053_)
);

INV_X4 _1364_ (
  .A(_1053_),
  .ZN(_1024_)
);

INV_X1 _1365_ (
  .A(_0987_),
  .ZN(_1027_)
);

INV_X1 _1366_ (
  .A(_0874_),
  .ZN(_0905_)
);

INV_X1 _1368_ (
  .A(_0785_),
  .ZN(_0786_)
);

INV_X1 _1370_ (
  .A(_0875_),
  .ZN(_0969_)
);

NAND2_X1 _1373_ (
  .A1(_0333_),
  .A2(_0358_),
  .ZN(_0822_)
);

INV_X1 _1374_ (
  .A(_0903_),
  .ZN(_0904_)
);

NAND2_X1 _1375_ (
  .A1(_0354_),
  .A2(_0358_),
  .ZN(_0920_)
);

INV_X1 _1376_ (
  .A(_0936_),
  .ZN(_0938_)
);

INV_X1 _1377_ (
  .A(_0968_),
  .ZN(_0970_)
);

INV_X1 _1378_ (
  .A(_1088_),
  .ZN(_0678_)
);

INV_X1 _1381_ (
  .A(_1152_),
  .ZN(_0787_)
);

INV_X1 _1382_ (
  .A(_1186_),
  .ZN(_0879_)
);

INV_X1 _1383_ (
  .A(_1193_),
  .ZN(_0916_)
);

NAND2_X1 _1384_ (
  .A1(_0356_),
  .A2(_0359_),
  .ZN(_1054_)
);

INV_X1 _1385_ (
  .A(_1029_),
  .ZN(_1067_)
);

INV_X1 _1386_ (
  .A(_0752_),
  .ZN(_0775_)
);

INV_X1 _1387_ (
  .A(_0769_),
  .ZN(_0771_)
);

INV_X1 _1388_ (
  .A(_0856_),
  .ZN(_0862_)
);

INV_X1 _1389_ (
  .A(_0884_),
  .ZN(_0890_)
);

INV_X1 _1390_ (
  .A(_0912_),
  .ZN(_0913_)
);

INV_X1 _1391_ (
  .A(_0950_),
  .ZN(_1204_)
);

INV_X1 _1392_ (
  .A(_0955_),
  .ZN(_0956_)
);

INV_X1 _1393_ (
  .A(_0985_),
  .ZN(_1211_)
);

INV_X1 _1394_ (
  .A(_0988_),
  .ZN(_0989_)
);

INV_X1 _1395_ (
  .A(_1026_),
  .ZN(_1028_)
);

INV_X1 _1396_ (
  .A(_1037_),
  .ZN(_1038_)
);

INV_X1 _1397_ (
  .A(_1056_),
  .ZN(_1057_)
);

INV_X1 _1398_ (
  .A(_1079_),
  .ZN(_1080_)
);

INV_X1 _1399_ (
  .A(_0689_),
  .ZN(_0699_)
);

INV_X1 _1400_ (
  .A(_0751_),
  .ZN(_0745_)
);

INV_X1 _1401_ (
  .A(_0776_),
  .ZN(_0770_)
);

INV_X1 _1402_ (
  .A(_0855_),
  .ZN(_0891_)
);

INV_X1 _1403_ (
  .A(_0883_),
  .ZN(_0924_)
);

INV_X1 _1404_ (
  .A(_0954_),
  .ZN(_0996_)
);

INV_X1 _1405_ (
  .A(_1007_),
  .ZN(_1039_)
);

INV_X1 _1406_ (
  .A(_1025_),
  .ZN(_1058_)
);

INV_X1 _1407_ (
  .A(_0702_),
  .ZN(_1141_)
);

INV_X1 _1408_ (
  .A(_0714_),
  .ZN(_0715_)
);

INV_X1 _1409_ (
  .A(_0711_),
  .ZN(_1150_)
);

INV_X1 _1410_ (
  .A(_0734_),
  .ZN(_1154_)
);

INV_X1 _1413_ (
  .A(_0723_),
  .ZN(_0774_)
);

INV_X1 _1414_ (
  .A(_0756_),
  .ZN(_0765_)
);

INV_X1 _1415_ (
  .A(_0728_),
  .ZN(_1163_)
);

INV_X1 _1416_ (
  .A(_0773_),
  .ZN(_0778_)
);

INV_X1 _1417_ (
  .A(_0789_),
  .ZN(_1171_)
);

INV_X1 _1418_ (
  .A(_0743_),
  .ZN(_0811_)
);

INV_X1 _1419_ (
  .A(_0820_),
  .ZN(_1179_)
);

INV_X1 _1420_ (
  .A(_0836_),
  .ZN(_0838_)
);

INV_X1 _1421_ (
  .A(_0809_),
  .ZN(_0837_)
);

INV_X1 _1422_ (
  .A(_0846_),
  .ZN(_0848_)
);

INV_X1 _1423_ (
  .A(_0869_),
  .ZN(_0908_)
);

INV_X1 _1424_ (
  .A(_0880_),
  .ZN(_1199_)
);

INV_X1 _1425_ (
  .A(_0946_),
  .ZN(_0947_)
);

INV_X1 _1426_ (
  .A(_0931_),
  .ZN(_0974_)
);

INV_X1 _1427_ (
  .A(_0945_),
  .ZN(_0982_)
);

INV_X1 _1428_ (
  .A(_0943_),
  .ZN(_1210_)
);

INV_X1 _1429_ (
  .A(_0991_),
  .ZN(_1216_)
);

INV_X1 _1430_ (
  .A(_0963_),
  .ZN(_1009_)
);

INV_X1 _1431_ (
  .A(_1017_),
  .ZN(_1018_)
);

INV_X1 _1432_ (
  .A(_0990_),
  .ZN(_1222_)
);

INV_X1 _1433_ (
  .A(_1046_),
  .ZN(_1047_)
);

INV_X1 _1434_ (
  .A(_1040_),
  .ZN(_1075_)
);

INV_X1 _1435_ (
  .A(_1082_),
  .ZN(_1083_)
);

INV_X1 _1436_ (
  .A(_0701_),
  .ZN(_0716_)
);

INV_X1 _1437_ (
  .A(_0762_),
  .ZN(_0766_)
);

INV_X1 _1438_ (
  .A(_0783_),
  .ZN(_0779_)
);

INV_X1 _1439_ (
  .A(_0788_),
  .ZN(_1165_)
);

INV_X1 _1440_ (
  .A(_0810_),
  .ZN(_0812_)
);

INV_X1 _1441_ (
  .A(_0761_),
  .ZN(_0813_)
);

INV_X1 _1442_ (
  .A(_0803_),
  .ZN(_0839_)
);

INV_X1 _1443_ (
  .A(_0819_),
  .ZN(_0849_)
);

INV_X1 _1444_ (
  .A(_0907_),
  .ZN(_0909_)
);

INV_X1 _1445_ (
  .A(_0914_),
  .ZN(_0948_)
);

INV_X1 _1446_ (
  .A(_0917_),
  .ZN(_1205_)
);

INV_X1 _1447_ (
  .A(_0935_),
  .ZN(_0973_)
);

INV_X1 _1448_ (
  .A(_0972_),
  .ZN(_0975_)
);

INV_X1 _1449_ (
  .A(_0939_),
  .ZN(_0976_)
);

INV_X1 _1450_ (
  .A(_0980_),
  .ZN(_0983_)
);

INV_X1 _1451_ (
  .A(_0967_),
  .ZN(_1006_)
);

INV_X1 _1452_ (
  .A(_0971_),
  .ZN(_1010_)
);

INV_X1 _1453_ (
  .A(_0902_),
  .ZN(_0942_)
);

INV_X1 _1454_ (
  .A(_1016_),
  .ZN(_1048_)
);

INV_X1 _1455_ (
  .A(_1045_),
  .ZN(_1084_)
);

INV_X1 _1456_ (
  .A(_1153_),
  .ZN(_0732_)
);

INV_X1 _1457_ (
  .A(_1170_),
  .ZN(_0790_)
);

INV_X1 _1458_ (
  .A(_1178_),
  .ZN(_0818_)
);

INV_X1 _1459_ (
  .A(_1187_),
  .ZN(_0844_)
);

INV_X1 _1460_ (
  .A(_1194_),
  .ZN(_0876_)
);

INV_X1 _1461_ (
  .A(_1219_),
  .ZN(_1015_)
);

INV_X1 _1462_ (
  .A(_1228_),
  .ZN(_1044_)
);

INV_X1 _1463_ (
  .A(_1140_),
  .ZN(_0700_)
);

INV_X1 _1464_ (
  .A(_1164_),
  .ZN(_0784_)
);

INV_X1 _1465_ (
  .A(_0941_),
  .ZN(_0937_)
);

INV_X1 _1466_ (
  .A(_1173_),
  .ZN(_0791_)
);

BUF_X1 _1467_ (
  .A(ena),
  .Z(_0367_)
);

BUF_X1 _1468_ (
  .A(_0367_),
  .Z(_0368_)
);

INV_X1 _1470_ (
  .A(\ext_mult_res[0] ),
  .ZN(_0370_)
);

BUF_X1 _1471_ (
  .A(_0367_),
  .Z(_0371_)
);

BUF_X1 _1472_ (
  .A(_0371_),
  .Z(_0372_)
);

BUF_X1 _1474_ (
  .A(_0367_),
  .Z(_0373_)
);

MUX2_X1 _1475_ (
  .A(\ext_mult_res[1] ),
  .B(_1133_),
  .S(_0373_),
  .Z(_0001_)
);

BUF_X4 _1476_ (
  .A(_0371_),
  .Z(_0374_)
);

NAND2_X1 _1477_ (
  .A1(_0374_),
  .A2(_1135_),
  .ZN(_0375_)
);

INV_X1 _1478_ (
  .A(\ext_mult_res[2] ),
  .ZN(_0376_)
);

OAI21_X1 _1479_ (
  .A(_0375_),
  .B1(_0376_),
  .B2(_0372_),
  .ZN(_0002_)
);

NAND2_X1 _1480_ (
  .A1(_0374_),
  .A2(_1137_),
  .ZN(_0377_)
);

INV_X1 _1481_ (
  .A(\ext_mult_res[3] ),
  .ZN(_0378_)
);

OAI21_X1 _1482_ (
  .A(_0377_),
  .B1(_0378_),
  .B2(_0372_),
  .ZN(_0003_)
);

NAND2_X1 _1483_ (
  .A1(_0374_),
  .A2(_1145_),
  .ZN(_0379_)
);

INV_X1 _1484_ (
  .A(\ext_mult_res[4] ),
  .ZN(_0380_)
);

OAI21_X1 _1485_ (
  .A(_0379_),
  .B1(_0380_),
  .B2(_0372_),
  .ZN(_0004_)
);

MUX2_X1 _1486_ (
  .A(\ext_mult_res[5] ),
  .B(_1149_),
  .S(_0373_),
  .Z(_0005_)
);

NAND2_X1 _1487_ (
  .A1(_0372_),
  .A2(_1160_),
  .ZN(_0381_)
);

INV_X1 _1488_ (
  .A(\ext_mult_res[6] ),
  .ZN(_0382_)
);

OAI21_X1 _1489_ (
  .A(_0381_),
  .B1(_0382_),
  .B2(_0372_),
  .ZN(_0006_)
);

NAND2_X1 _1490_ (
  .A1(_0374_),
  .A2(_1234_),
  .ZN(_0383_)
);

INV_X1 _1491_ (
  .A(\ext_mult_res[7] ),
  .ZN(_0384_)
);

OAI21_X1 _1492_ (
  .A(_0383_),
  .B1(_0384_),
  .B2(_0372_),
  .ZN(_0007_)
);

INV_X1 _1493_ (
  .A(_0367_),
  .ZN(_0385_)
);

NAND2_X1 _1494_ (
  .A1(_0385_),
  .A2(\ext_mult_res[8] ),
  .ZN(_0386_)
);

BUF_X1 _1495_ (
  .A(_0385_),
  .Z(_0387_)
);

OAI21_X1 _1496_ (
  .A(_0386_),
  .B1(_0794_),
  .B2(_0387_),
  .ZN(_0008_)
);

INV_X1 _1497_ (
  .A(_0793_),
  .ZN(_0388_)
);

NAND2_X1 _1498_ (
  .A1(_0388_),
  .A2(_1185_),
  .ZN(_0389_)
);

INV_X1 _1499_ (
  .A(_1185_),
  .ZN(_0390_)
);

NAND2_X1 _1500_ (
  .A1(_0390_),
  .A2(_0793_),
  .ZN(_0391_)
);

NAND3_X1 _1501_ (
  .A1(_0389_),
  .A2(_0391_),
  .A3(_0374_),
  .ZN(_0392_)
);

INV_X1 _1502_ (
  .A(\ext_mult_res[9] ),
  .ZN(_0393_)
);

OAI21_X1 _1503_ (
  .A(_0392_),
  .B1(_0393_),
  .B2(_0372_),
  .ZN(_0009_)
);

NOR2_X1 _1504_ (
  .A1(\ext_mult_res[10] ),
  .A2(_0373_),
  .ZN(_0394_)
);

INV_X1 _1505_ (
  .A(_1184_),
  .ZN(_0395_)
);

INV_X1 _1506_ (
  .A(_1174_),
  .ZN(_0396_)
);

OAI21_X1 _1507_ (
  .A(_0395_),
  .B1(_0390_),
  .B2(_0396_),
  .ZN(_0397_)
);

INV_X1 _1508_ (
  .A(_0397_),
  .ZN(_0398_)
);

NAND2_X1 _1509_ (
  .A1(_1185_),
  .A2(_1175_),
  .ZN(_0399_)
);

OAI21_X1 _1510_ (
  .A(_0398_),
  .B1(_0792_),
  .B2(_0399_),
  .ZN(_0400_)
);

BUF_X1 _1511_ (
  .A(_1191_),
  .Z(_0401_)
);

XNOR2_X1 _1512_ (
  .A(_0400_),
  .B(_0401_),
  .ZN(_0402_)
);

BUF_X1 _1513_ (
  .A(_0371_),
  .Z(_0403_)
);

AOI21_X1 _1514_ (
  .A(_0394_),
  .B1(_0402_),
  .B2(_0403_),
  .ZN(_0010_)
);

NOR2_X1 _1515_ (
  .A1(\ext_mult_res[11] ),
  .A2(_0373_),
  .ZN(_0404_)
);

INV_X1 _1516_ (
  .A(_1190_),
  .ZN(_0405_)
);

INV_X1 _1517_ (
  .A(_0401_),
  .ZN(_0406_)
);

OAI21_X1 _1518_ (
  .A(_0405_),
  .B1(_0406_),
  .B2(_0395_),
  .ZN(_0407_)
);

NAND2_X1 _1519_ (
  .A1(_1185_),
  .A2(_0401_),
  .ZN(_0408_)
);

INV_X1 _1520_ (
  .A(_0408_),
  .ZN(_0409_)
);

AOI21_X1 _1521_ (
  .A(_0407_),
  .B1(_0409_),
  .B2(_0388_),
  .ZN(_0410_)
);

INV_X1 _1522_ (
  .A(_1198_),
  .ZN(_0411_)
);

XNOR2_X1 _1523_ (
  .A(_0410_),
  .B(_0411_),
  .ZN(_0412_)
);

AOI21_X1 _1524_ (
  .A(_0404_),
  .B1(_0412_),
  .B2(_0403_),
  .ZN(_0011_)
);

NOR2_X1 _1525_ (
  .A1(\ext_mult_res[12] ),
  .A2(_0373_),
  .ZN(_0413_)
);

INV_X1 _1526_ (
  .A(_1197_),
  .ZN(_0414_)
);

OAI21_X1 _1527_ (
  .A(_0414_),
  .B1(_0411_),
  .B2(_0405_),
  .ZN(_0415_)
);

INV_X1 _1528_ (
  .A(_0415_),
  .ZN(_0416_)
);

NAND2_X1 _1529_ (
  .A1(_0401_),
  .A2(_1198_),
  .ZN(_0417_)
);

OAI21_X1 _1530_ (
  .A(_0416_),
  .B1(_0398_),
  .B2(_0417_),
  .ZN(_0418_)
);

NOR2_X1 _1531_ (
  .A1(_0399_),
  .A2(_0417_),
  .ZN(_0419_)
);

AOI21_X1 _1532_ (
  .A(_0418_),
  .B1(_0419_),
  .B2(_1177_),
  .ZN(_0420_)
);

INV_X1 _1533_ (
  .A(_1203_),
  .ZN(_0421_)
);

XNOR2_X1 _1534_ (
  .A(_0420_),
  .B(_0421_),
  .ZN(_0422_)
);

AOI21_X1 _1535_ (
  .A(_0413_),
  .B1(_0422_),
  .B2(_0403_),
  .ZN(_0012_)
);

NOR2_X1 _1536_ (
  .A1(\ext_mult_res[13] ),
  .A2(_0373_),
  .ZN(_0423_)
);

INV_X1 _1537_ (
  .A(_1202_),
  .ZN(_0424_)
);

OAI21_X1 _1538_ (
  .A(_0424_),
  .B1(_0421_),
  .B2(_0414_),
  .ZN(_0425_)
);

INV_X1 _1539_ (
  .A(_0425_),
  .ZN(_0426_)
);

INV_X1 _1540_ (
  .A(_0407_),
  .ZN(_0427_)
);

NAND2_X1 _1541_ (
  .A1(_1198_),
  .A2(_1203_),
  .ZN(_0428_)
);

OAI21_X1 _1542_ (
  .A(_0426_),
  .B1(_0427_),
  .B2(_0428_),
  .ZN(_0429_)
);

NOR2_X1 _1543_ (
  .A1(_0408_),
  .A2(_0428_),
  .ZN(_0430_)
);

AOI21_X1 _1544_ (
  .A(_0429_),
  .B1(_0430_),
  .B2(_0388_),
  .ZN(_0431_)
);

INV_X1 _1545_ (
  .A(_1209_),
  .ZN(_0432_)
);

XNOR2_X1 _1546_ (
  .A(_0431_),
  .B(_0432_),
  .ZN(_0433_)
);

AOI21_X1 _1547_ (
  .A(_0423_),
  .B1(_0433_),
  .B2(_0403_),
  .ZN(_0013_)
);

NOR2_X1 _1548_ (
  .A1(\ext_mult_res[14] ),
  .A2(_0373_),
  .ZN(_0434_)
);

INV_X1 _1549_ (
  .A(_1208_),
  .ZN(_0435_)
);

OAI21_X1 _1550_ (
  .A(_0435_),
  .B1(_0432_),
  .B2(_0424_),
  .ZN(_0436_)
);

INV_X1 _1551_ (
  .A(_0436_),
  .ZN(_0437_)
);

NAND2_X1 _1552_ (
  .A1(_1203_),
  .A2(_1209_),
  .ZN(_0438_)
);

OAI21_X1 _1553_ (
  .A(_0437_),
  .B1(_0416_),
  .B2(_0438_),
  .ZN(_0439_)
);

NOR2_X1 _1554_ (
  .A1(_0417_),
  .A2(_0438_),
  .ZN(_0440_)
);

AOI21_X1 _1555_ (
  .A(_0439_),
  .B1(_0440_),
  .B2(_0400_),
  .ZN(_0441_)
);

INV_X1 _1556_ (
  .A(_1215_),
  .ZN(_0442_)
);

XNOR2_X1 _1557_ (
  .A(_0441_),
  .B(_0442_),
  .ZN(_0443_)
);

AOI21_X1 _1558_ (
  .A(_0434_),
  .B1(_0443_),
  .B2(_0403_),
  .ZN(_0014_)
);

NAND2_X1 _1559_ (
  .A1(_1209_),
  .A2(_1215_),
  .ZN(_0444_)
);

NOR3_X1 _1560_ (
  .A1(_0410_),
  .A2(_0428_),
  .A3(_0444_),
  .ZN(_0445_)
);

INV_X1 _1561_ (
  .A(_1214_),
  .ZN(_0446_)
);

OAI21_X1 _1562_ (
  .A(_0446_),
  .B1(_0442_),
  .B2(_0435_),
  .ZN(_0447_)
);

INV_X1 _1563_ (
  .A(_0447_),
  .ZN(_0448_)
);

OAI21_X1 _1564_ (
  .A(_0448_),
  .B1(_0426_),
  .B2(_0444_),
  .ZN(_0449_)
);

OR2_X1 _1565_ (
  .A1(_0445_),
  .A2(_0449_),
  .ZN(_0450_)
);

BUF_X1 _1566_ (
  .A(_1221_),
  .Z(_0451_)
);

OR2_X1 _1567_ (
  .A1(_0450_),
  .A2(_0451_),
  .ZN(_0452_)
);

NAND2_X1 _1568_ (
  .A1(_0450_),
  .A2(_0451_),
  .ZN(_0453_)
);

NAND3_X1 _1569_ (
  .A1(_0452_),
  .A2(_0374_),
  .A3(_0453_),
  .ZN(_0454_)
);

INV_X1 _1570_ (
  .A(\ext_mult_res[15] ),
  .ZN(_0455_)
);

OAI21_X1 _1571_ (
  .A(_0454_),
  .B1(_0455_),
  .B2(_0372_),
  .ZN(_0015_)
);

NOR2_X1 _1572_ (
  .A1(\ext_mult_res[16] ),
  .A2(_0373_),
  .ZN(_0456_)
);

INV_X1 _1573_ (
  .A(_1220_),
  .ZN(_0457_)
);

INV_X1 _1574_ (
  .A(_0451_),
  .ZN(_0458_)
);

OAI21_X1 _1575_ (
  .A(_0457_),
  .B1(_0458_),
  .B2(_0446_),
  .ZN(_0459_)
);

INV_X1 _1576_ (
  .A(_0459_),
  .ZN(_0460_)
);

NAND2_X1 _1577_ (
  .A1(_1215_),
  .A2(_0451_),
  .ZN(_0461_)
);

OAI21_X1 _1578_ (
  .A(_0460_),
  .B1(_0437_),
  .B2(_0461_),
  .ZN(_0462_)
);

NOR2_X1 _1579_ (
  .A1(_0438_),
  .A2(_0461_),
  .ZN(_0463_)
);

AOI21_X1 _1580_ (
  .A(_0462_),
  .B1(_0463_),
  .B2(_0418_),
  .ZN(_0464_)
);

NAND3_X1 _1581_ (
  .A1(_0419_),
  .A2(_0463_),
  .A3(_1177_),
  .ZN(_0465_)
);

NAND2_X1 _1582_ (
  .A1(_0464_),
  .A2(_0465_),
  .ZN(_0466_)
);

BUF_X1 _1583_ (
  .A(_1230_),
  .Z(_0467_)
);

XNOR2_X1 _1584_ (
  .A(_0466_),
  .B(_0467_),
  .ZN(_0468_)
);

AOI21_X1 _1585_ (
  .A(_0456_),
  .B1(_0468_),
  .B2(_0403_),
  .ZN(_0016_)
);

NOR2_X1 _1586_ (
  .A1(\ext_mult_res[17] ),
  .A2(_0373_),
  .ZN(_0469_)
);

INV_X1 _1587_ (
  .A(_1229_),
  .ZN(_0470_)
);

INV_X1 _1588_ (
  .A(_0467_),
  .ZN(_0471_)
);

NAND2_X1 _1589_ (
  .A1(_0451_),
  .A2(_0467_),
  .ZN(_0472_)
);

OAI221_X1 _1590_ (
  .A(_0470_),
  .B1(_0457_),
  .B2(_0471_),
  .C1(_0448_),
  .C2(_0472_),
  .ZN(_0473_)
);

INV_X1 _1591_ (
  .A(_0473_),
  .ZN(_0474_)
);

NOR2_X1 _1592_ (
  .A1(_0444_),
  .A2(_0472_),
  .ZN(_0475_)
);

NAND2_X1 _1593_ (
  .A1(_0429_),
  .A2(_0475_),
  .ZN(_0476_)
);

NAND3_X1 _1594_ (
  .A1(_0430_),
  .A2(_0475_),
  .A3(_0388_),
  .ZN(_0477_)
);

NAND3_X1 _1595_ (
  .A1(_0474_),
  .A2(_0476_),
  .A3(_0477_),
  .ZN(_0478_)
);

BUF_X1 _1596_ (
  .A(_1233_),
  .Z(_0479_)
);

XNOR2_X1 _1597_ (
  .A(_0478_),
  .B(_0479_),
  .ZN(_0480_)
);

AOI21_X1 _1598_ (
  .A(_0469_),
  .B1(_0480_),
  .B2(_0403_),
  .ZN(_0017_)
);

INV_X1 _1599_ (
  .A(_1061_),
  .ZN(_0481_)
);

INV_X1 _1600_ (
  .A(_1070_),
  .ZN(_0482_)
);

NAND2_X1 _1601_ (
  .A1(_0481_),
  .A2(_0482_),
  .ZN(_0483_)
);

NAND2_X1 _1602_ (
  .A1(_1061_),
  .A2(_1070_),
  .ZN(_0484_)
);

NAND2_X1 _1603_ (
  .A1(_0483_),
  .A2(_0484_),
  .ZN(_0485_)
);

INV_X1 _1604_ (
  .A(_0485_),
  .ZN(_0486_)
);

INV_X1 _1605_ (
  .A(_1081_),
  .ZN(_0487_)
);

NAND2_X1 _1606_ (
  .A1(_0487_),
  .A2(_1055_),
  .ZN(_0488_)
);

INV_X1 _1607_ (
  .A(_1055_),
  .ZN(_0489_)
);

NAND2_X1 _1608_ (
  .A1(_0489_),
  .A2(_1081_),
  .ZN(_0490_)
);

NAND2_X1 _1609_ (
  .A1(_0488_),
  .A2(_0490_),
  .ZN(_0491_)
);

NAND2_X1 _1610_ (
  .A1(_0486_),
  .A2(_0491_),
  .ZN(_0492_)
);

XNOR2_X1 _1611_ (
  .A(_1081_),
  .B(_1055_),
  .ZN(_0493_)
);

NAND2_X1 _1612_ (
  .A1(_0493_),
  .A2(_0485_),
  .ZN(_0494_)
);

NAND2_X1 _1613_ (
  .A1(_0492_),
  .A2(_0494_),
  .ZN(_0495_)
);

INV_X1 _1614_ (
  .A(_1224_),
  .ZN(_0496_)
);

NAND2_X1 _1615_ (
  .A1(_0496_),
  .A2(_1027_),
  .ZN(_0497_)
);

NAND2_X1 _1616_ (
  .A1(_1224_),
  .A2(_0987_),
  .ZN(_0498_)
);

NAND2_X1 _1617_ (
  .A1(_0497_),
  .A2(_0498_),
  .ZN(_0499_)
);

NAND2_X1 _1618_ (
  .A1(_0499_),
  .A2(_1023_),
  .ZN(_0500_)
);

NAND3_X1 _1619_ (
  .A1(_0497_),
  .A2(_1052_),
  .A3(_0498_),
  .ZN(_0501_)
);

NAND2_X2 _1620_ (
  .A1(_0500_),
  .A2(_0501_),
  .ZN(_0502_)
);

XNOR2_X1 _1621_ (
  .A(_0495_),
  .B(_0502_),
  .ZN(_0503_)
);

INV_X1 _1622_ (
  .A(_1005_),
  .ZN(_0504_)
);

XNOR2_X1 _1623_ (
  .A(_0504_),
  .B(_1059_),
  .ZN(_0505_)
);

XNOR2_X1 _1624_ (
  .A(_1063_),
  .B(_1065_),
  .ZN(_0506_)
);

NAND2_X1 _1625_ (
  .A1(_0505_),
  .A2(_0506_),
  .ZN(_0507_)
);

NAND2_X1 _1626_ (
  .A1(_1063_),
  .A2(_1065_),
  .ZN(_0508_)
);

INV_X1 _1627_ (
  .A(_0508_),
  .ZN(_0509_)
);

NOR2_X1 _1628_ (
  .A1(_1063_),
  .A2(_1065_),
  .ZN(_0510_)
);

NOR2_X1 _1629_ (
  .A1(_0509_),
  .A2(_0510_),
  .ZN(_0511_)
);

XNOR2_X1 _1630_ (
  .A(_1005_),
  .B(_1059_),
  .ZN(_0512_)
);

NAND2_X1 _1631_ (
  .A1(_0511_),
  .A2(_0512_),
  .ZN(_0513_)
);

NAND2_X1 _1632_ (
  .A1(_0507_),
  .A2(_0513_),
  .ZN(_0514_)
);

INV_X1 _1633_ (
  .A(_0514_),
  .ZN(_0515_)
);

NAND2_X2 _1637_ (
  .A1(_0518_),
  .A2(_1053_),
  .ZN(_0519_)
);

NAND2_X2 _1639_ (
  .A1(_0519_),
  .A2(_0520_),
  .ZN(_0521_)
);

NAND2_X1 _1640_ (
  .A1(_0515_),
  .A2(_0521_),
  .ZN(_0522_)
);

NAND2_X2 _1641_ (
  .A1(_0518_),
  .A2(_1024_),
  .ZN(_0523_)
);

INV_X1 _1642_ (
  .A(_0358_),
  .ZN(_0524_)
);

NAND2_X2 _1644_ (
  .A1(_0523_),
  .A2(_0525_),
  .ZN(_0526_)
);

NAND2_X1 _1645_ (
  .A1(_0526_),
  .A2(_0514_),
  .ZN(_0527_)
);

NAND2_X2 _1646_ (
  .A1(_0522_),
  .A2(_0527_),
  .ZN(_0528_)
);

NAND2_X1 _1647_ (
  .A1(_0503_),
  .A2(_0528_),
  .ZN(_0529_)
);

NAND2_X1 _1648_ (
  .A1(_0515_),
  .A2(_0526_),
  .ZN(_0530_)
);

NAND2_X1 _1649_ (
  .A1(_0521_),
  .A2(_0514_),
  .ZN(_0531_)
);

NAND2_X2 _1650_ (
  .A1(_0530_),
  .A2(_0531_),
  .ZN(_0532_)
);

XNOR2_X1 _1651_ (
  .A(_0491_),
  .B(_0485_),
  .ZN(_0533_)
);

NAND2_X1 _1652_ (
  .A1(_0533_),
  .A2(_0502_),
  .ZN(_0534_)
);

INV_X1 _1653_ (
  .A(_0502_),
  .ZN(_0535_)
);

NAND2_X1 _1654_ (
  .A1(_0495_),
  .A2(_0535_),
  .ZN(_0536_)
);

NAND2_X1 _1655_ (
  .A1(_0534_),
  .A2(_0536_),
  .ZN(_0537_)
);

NAND2_X1 _1656_ (
  .A1(_0532_),
  .A2(_0537_),
  .ZN(_0538_)
);

NAND2_X1 _1657_ (
  .A1(_0529_),
  .A2(_0538_),
  .ZN(_0539_)
);

OR2_X1 _1658_ (
  .A1(_1086_),
  .A2(_1078_),
  .ZN(_0540_)
);

NAND2_X1 _1659_ (
  .A1(_1078_),
  .A2(_1086_),
  .ZN(_0541_)
);

XOR2_X1 _1664_ (
  .A(_1068_),
  .B(_1231_),
  .Z(_0546_)
);

INV_X1 _1665_ (
  .A(_0546_),
  .ZN(_0547_)
);

NAND2_X2 _1666_ (
  .A1(_0545_),
  .A2(_0547_),
  .ZN(_0548_)
);

NAND2_X2 _1668_ (
  .A1(_0548_),
  .A2(_0549_),
  .ZN(_0550_)
);

XNOR2_X1 _1669_ (
  .A(_0967_),
  .B(_0903_),
  .ZN(_0551_)
);

XNOR2_X1 _1670_ (
  .A(_0874_),
  .B(_1073_),
  .ZN(_0552_)
);

XNOR2_X1 _1671_ (
  .A(_0551_),
  .B(_0552_),
  .ZN(_0553_)
);

INV_X1 _1672_ (
  .A(_0553_),
  .ZN(_0554_)
);

NAND2_X2 _1673_ (
  .A1(_0550_),
  .A2(_0554_),
  .ZN(_0555_)
);

NAND3_X1 _1674_ (
  .A1(_0548_),
  .A2(_0549_),
  .A3(_0553_),
  .ZN(_0556_)
);

NAND2_X2 _1675_ (
  .A1(_0555_),
  .A2(_0556_),
  .ZN(_0557_)
);

INV_X1 _1676_ (
  .A(_0557_),
  .ZN(_0558_)
);

NAND2_X2 _1677_ (
  .A1(_0539_),
  .A2(_0558_),
  .ZN(_0559_)
);

NAND2_X1 _1678_ (
  .A1(_0503_),
  .A2(_0532_),
  .ZN(_0560_)
);

NAND2_X1 _1679_ (
  .A1(_0528_),
  .A2(_0537_),
  .ZN(_0561_)
);

NAND2_X2 _1680_ (
  .A1(_0560_),
  .A2(_0561_),
  .ZN(_0562_)
);

NAND2_X2 _1681_ (
  .A1(_0562_),
  .A2(_0557_),
  .ZN(_0563_)
);

NAND2_X2 _1682_ (
  .A1(_0559_),
  .A2(_0563_),
  .ZN(_0564_)
);

INV_X1 _1683_ (
  .A(_0479_),
  .ZN(_0565_)
);

NOR3_X1 _1684_ (
  .A1(_0461_),
  .A2(_0471_),
  .A3(_0565_),
  .ZN(_0566_)
);

NAND3_X1 _1685_ (
  .A1(_0400_),
  .A2(_0440_),
  .A3(_0566_),
  .ZN(_0567_)
);

NAND3_X1 _1686_ (
  .A1(_0459_),
  .A2(_0467_),
  .A3(_0479_),
  .ZN(_0568_)
);

INV_X1 _1687_ (
  .A(_1232_),
  .ZN(_0569_)
);

NAND2_X1 _1688_ (
  .A1(_0479_),
  .A2(_1229_),
  .ZN(_0570_)
);

NAND3_X1 _1689_ (
  .A1(_0568_),
  .A2(_0569_),
  .A3(_0570_),
  .ZN(_0571_)
);

INV_X1 _1690_ (
  .A(_0571_),
  .ZN(_0572_)
);

NAND2_X1 _1691_ (
  .A1(_0439_),
  .A2(_0566_),
  .ZN(_0573_)
);

AND3_X1 _1692_ (
  .A1(_0567_),
  .A2(_0572_),
  .A3(_0573_),
  .ZN(_0574_)
);

INV_X1 _1693_ (
  .A(_0574_),
  .ZN(_0575_)
);

NAND2_X2 _1694_ (
  .A1(_0564_),
  .A2(_0575_),
  .ZN(_0576_)
);

NAND3_X1 _1695_ (
  .A1(_0559_),
  .A2(_0563_),
  .A3(_0574_),
  .ZN(_0577_)
);

NAND3_X1 _1696_ (
  .A1(_0576_),
  .A2(_0577_),
  .A3(_0374_),
  .ZN(_0578_)
);

NAND2_X1 _1697_ (
  .A1(_0387_),
  .A2(\ext_mult_res[18] ),
  .ZN(_0579_)
);

NAND2_X1 _1698_ (
  .A1(_0578_),
  .A2(_0579_),
  .ZN(_0018_)
);

NAND2_X1 _1699_ (
  .A1(_0385_),
  .A2(result[0]),
  .ZN(_0580_)
);

BUF_X1 _1700_ (
  .A(dclr),
  .Z(_0581_)
);

OAI21_X1 _1701_ (
  .A(_0368_),
  .B1(_1089_),
  .B2(_0581_),
  .ZN(_0582_)
);

INV_X1 _1702_ (
  .A(_0581_),
  .ZN(_0583_)
);

BUF_X1 _1703_ (
  .A(_0583_),
  .Z(_0584_)
);

NOR2_X1 _1704_ (
  .A1(_0584_),
  .A2(\ext_mult_res[0] ),
  .ZN(_0585_)
);

OAI21_X1 _1705_ (
  .A(_0580_),
  .B1(_0582_),
  .B2(_0585_),
  .ZN(_0019_)
);

NAND2_X1 _1706_ (
  .A1(_0385_),
  .A2(result[1]),
  .ZN(_0586_)
);

OAI21_X1 _1707_ (
  .A(_0368_),
  .B1(_0581_),
  .B2(_0680_),
  .ZN(_0587_)
);

NOR2_X1 _1708_ (
  .A1(_0584_),
  .A2(\ext_mult_res[1] ),
  .ZN(_0588_)
);

OAI21_X1 _1709_ (
  .A(_0586_),
  .B1(_0587_),
  .B2(_0588_),
  .ZN(_0020_)
);

INV_X1 _1710_ (
  .A(_1093_),
  .ZN(_0589_)
);

NOR2_X1 _1711_ (
  .A1(_0589_),
  .A2(_0679_),
  .ZN(_0590_)
);

INV_X1 _1712_ (
  .A(_0590_),
  .ZN(_0591_)
);

NAND2_X1 _1713_ (
  .A1(_0589_),
  .A2(_0679_),
  .ZN(_0592_)
);

NAND3_X1 _1714_ (
  .A1(_0591_),
  .A2(_0583_),
  .A3(_0592_),
  .ZN(_0593_)
);

BUF_X2 _1715_ (
  .A(_0583_),
  .Z(_0594_)
);

OAI21_X1 _1716_ (
  .A(_0593_),
  .B1(_0594_),
  .B2(_0376_),
  .ZN(_0595_)
);

MUX2_X1 _1717_ (
  .A(result[2]),
  .B(_0595_),
  .S(_0373_),
  .Z(_0021_)
);

OAI21_X1 _1718_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(_0378_),
  .ZN(_0596_)
);

NAND2_X1 _1719_ (
  .A1(_1088_),
  .A2(_1091_),
  .ZN(_0597_)
);

INV_X1 _1720_ (
  .A(_1090_),
  .ZN(_0598_)
);

INV_X1 _1721_ (
  .A(_1092_),
  .ZN(_0599_)
);

NAND3_X1 _1722_ (
  .A1(_0597_),
  .A2(_0598_),
  .A3(_0599_),
  .ZN(_0600_)
);

NAND2_X1 _1723_ (
  .A1(_0589_),
  .A2(_0599_),
  .ZN(_0601_)
);

NAND2_X1 _1724_ (
  .A1(_0600_),
  .A2(_0601_),
  .ZN(_0602_)
);

XNOR2_X1 _1725_ (
  .A(_0602_),
  .B(_1095_),
  .ZN(_0603_)
);

BUF_X1 _1726_ (
  .A(_0583_),
  .Z(_0604_)
);

AOI21_X1 _1727_ (
  .A(_0596_),
  .B1(_0603_),
  .B2(_0604_),
  .ZN(_0605_)
);

INV_X1 _1728_ (
  .A(result[3]),
  .ZN(_0606_)
);

AOI21_X1 _1729_ (
  .A(_0605_),
  .B1(_0606_),
  .B2(_0387_),
  .ZN(_0022_)
);

OAI21_X1 _1730_ (
  .A(_0367_),
  .B1(_0583_),
  .B2(_0380_),
  .ZN(_0607_)
);

INV_X1 _1731_ (
  .A(_1094_),
  .ZN(_0608_)
);

INV_X1 _1732_ (
  .A(_1095_),
  .ZN(_0609_)
);

OAI21_X1 _1733_ (
  .A(_0608_),
  .B1(_0609_),
  .B2(_0599_),
  .ZN(_0610_)
);

INV_X1 _1734_ (
  .A(_0610_),
  .ZN(_0611_)
);

OAI21_X4 _1735_ (
  .A(_0611_),
  .B1(_0609_),
  .B2(_0591_),
  .ZN(_0612_)
);

INV_X1 _1736_ (
  .A(_1097_),
  .ZN(_0613_)
);

XNOR2_X1 _1737_ (
  .A(_0612_),
  .B(_0613_),
  .ZN(_0614_)
);

AOI21_X1 _1738_ (
  .A(_0607_),
  .B1(_0614_),
  .B2(_0604_),
  .ZN(_0615_)
);

INV_X1 _1739_ (
  .A(result[4]),
  .ZN(_0616_)
);

AOI21_X1 _1740_ (
  .A(_0615_),
  .B1(_0616_),
  .B2(_0387_),
  .ZN(_0023_)
);

NAND2_X1 _1741_ (
  .A1(_1095_),
  .A2(_1097_),
  .ZN(_0617_)
);

INV_X1 _1742_ (
  .A(_0617_),
  .ZN(_0618_)
);

NAND3_X1 _1743_ (
  .A1(_0600_),
  .A2(_0601_),
  .A3(_0618_),
  .ZN(_0619_)
);

INV_X1 _1744_ (
  .A(_1096_),
  .ZN(_0620_)
);

OAI21_X1 _1745_ (
  .A(_0620_),
  .B1(_0613_),
  .B2(_0608_),
  .ZN(_0621_)
);

INV_X1 _1746_ (
  .A(_0621_),
  .ZN(_0622_)
);

NAND2_X1 _1747_ (
  .A1(_0619_),
  .A2(_0622_),
  .ZN(_0623_)
);

BUF_X2 _1748_ (
  .A(_1099_),
  .Z(_0624_)
);

XNOR2_X1 _1749_ (
  .A(_0623_),
  .B(_0624_),
  .ZN(_0625_)
);

AOI21_X1 _1750_ (
  .A(_0385_),
  .B1(_0625_),
  .B2(_0594_),
  .ZN(_0626_)
);

OAI21_X1 _1751_ (
  .A(_0626_),
  .B1(_0584_),
  .B2(\ext_mult_res[5] ),
  .ZN(_0627_)
);

INV_X1 _1752_ (
  .A(result[5]),
  .ZN(_0628_)
);

OAI21_X1 _1753_ (
  .A(_0627_),
  .B1(_0403_),
  .B2(_0628_),
  .ZN(_0024_)
);

INV_X1 _1754_ (
  .A(_1098_),
  .ZN(_0629_)
);

INV_X1 _1755_ (
  .A(_0624_),
  .ZN(_0630_)
);

OAI21_X1 _1756_ (
  .A(_0629_),
  .B1(_0630_),
  .B2(_0620_),
  .ZN(_0631_)
);

INV_X1 _1757_ (
  .A(_0631_),
  .ZN(_0632_)
);

INV_X1 _1758_ (
  .A(_0612_),
  .ZN(_0633_)
);

NAND2_X1 _1759_ (
  .A1(_1097_),
  .A2(_0624_),
  .ZN(_0634_)
);

OAI21_X1 _1760_ (
  .A(_0632_),
  .B1(_0633_),
  .B2(_0634_),
  .ZN(_0635_)
);

CLKBUF_X2 _1761_ (
  .A(_1101_),
  .Z(_0636_)
);

XNOR2_X1 _1762_ (
  .A(_0635_),
  .B(_0636_),
  .ZN(_0041_)
);

NAND2_X1 _1763_ (
  .A1(_0041_),
  .A2(_0604_),
  .ZN(_0042_)
);

NAND2_X1 _1764_ (
  .A1(_0382_),
  .A2(_0581_),
  .ZN(_0043_)
);

NAND3_X1 _1765_ (
  .A1(_0042_),
  .A2(_0374_),
  .A3(_0043_),
  .ZN(_0044_)
);

INV_X1 _1766_ (
  .A(result[6]),
  .ZN(_0045_)
);

OAI21_X1 _1767_ (
  .A(_0044_),
  .B1(_0403_),
  .B2(_0045_),
  .ZN(_0025_)
);

NAND2_X1 _1768_ (
  .A1(_0636_),
  .A2(_1098_),
  .ZN(_0046_)
);

INV_X1 _1769_ (
  .A(_1100_),
  .ZN(_0047_)
);

NAND2_X1 _1770_ (
  .A1(_0046_),
  .A2(_0047_),
  .ZN(_0048_)
);

INV_X1 _1771_ (
  .A(_0048_),
  .ZN(_0049_)
);

NAND2_X1 _1772_ (
  .A1(_0624_),
  .A2(_0636_),
  .ZN(_0050_)
);

OAI21_X1 _1773_ (
  .A(_0049_),
  .B1(_0622_),
  .B2(_0050_),
  .ZN(_0051_)
);

INV_X1 _1774_ (
  .A(_0051_),
  .ZN(_0052_)
);

OAI21_X1 _1775_ (
  .A(_0052_),
  .B1(_0619_),
  .B2(_0050_),
  .ZN(_0053_)
);

BUF_X2 _1776_ (
  .A(_1103_),
  .Z(_0054_)
);

XNOR2_X1 _1777_ (
  .A(_0053_),
  .B(_0054_),
  .ZN(_0055_)
);

NAND2_X1 _1778_ (
  .A1(_0055_),
  .A2(_0604_),
  .ZN(_0056_)
);

NAND2_X1 _1779_ (
  .A1(_0384_),
  .A2(_0581_),
  .ZN(_0057_)
);

NAND3_X1 _1780_ (
  .A1(_0056_),
  .A2(_0374_),
  .A3(_0057_),
  .ZN(_0058_)
);

INV_X1 _1781_ (
  .A(result[7]),
  .ZN(_0059_)
);

OAI21_X1 _1782_ (
  .A(_0058_),
  .B1(_0403_),
  .B2(_0059_),
  .ZN(_0026_)
);

NAND2_X1 _1783_ (
  .A1(_0385_),
  .A2(result[8]),
  .ZN(_0060_)
);

INV_X1 _1784_ (
  .A(_1102_),
  .ZN(_0061_)
);

INV_X1 _1785_ (
  .A(_0054_),
  .ZN(_0062_)
);

OAI21_X1 _1786_ (
  .A(_0061_),
  .B1(_0062_),
  .B2(_0047_),
  .ZN(_0063_)
);

INV_X1 _1787_ (
  .A(_0063_),
  .ZN(_0064_)
);

NAND2_X1 _1788_ (
  .A1(_0636_),
  .A2(_0054_),
  .ZN(_0065_)
);

OAI21_X1 _1789_ (
  .A(_0064_),
  .B1(_0632_),
  .B2(_0065_),
  .ZN(_0066_)
);

INV_X1 _1790_ (
  .A(_0066_),
  .ZN(_0067_)
);

NOR2_X1 _1791_ (
  .A1(_0634_),
  .A2(_0065_),
  .ZN(_0068_)
);

INV_X1 _1792_ (
  .A(_0068_),
  .ZN(_0069_)
);

OAI21_X1 _1793_ (
  .A(_0067_),
  .B1(_0633_),
  .B2(_0069_),
  .ZN(_0070_)
);

INV_X1 _1794_ (
  .A(_1105_),
  .ZN(_0071_)
);

XNOR2_X1 _1795_ (
  .A(_0070_),
  .B(_0071_),
  .ZN(_0072_)
);

OAI21_X1 _1796_ (
  .A(_0368_),
  .B1(_0072_),
  .B2(_0581_),
  .ZN(_0073_)
);

NOR2_X1 _1797_ (
  .A1(_0584_),
  .A2(\ext_mult_res[8] ),
  .ZN(_0074_)
);

OAI21_X1 _1798_ (
  .A(_0060_),
  .B1(_0073_),
  .B2(_0074_),
  .ZN(_0027_)
);

OAI21_X1 _1799_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[9] ),
  .ZN(_0075_)
);

INV_X1 _1800_ (
  .A(_0075_),
  .ZN(_0076_)
);

NAND2_X2 _1801_ (
  .A1(_0054_),
  .A2(_1105_),
  .ZN(_0077_)
);

INV_X1 _1802_ (
  .A(_0077_),
  .ZN(_0078_)
);

NAND2_X1 _1803_ (
  .A1(_0053_),
  .A2(_0078_),
  .ZN(_0079_)
);

INV_X1 _1804_ (
  .A(_1104_),
  .ZN(_0080_)
);

OAI21_X1 _1805_ (
  .A(_0080_),
  .B1(_0071_),
  .B2(_0061_),
  .ZN(_0081_)
);

INV_X1 _1806_ (
  .A(_0081_),
  .ZN(_0082_)
);

NAND2_X1 _1807_ (
  .A1(_0079_),
  .A2(_0082_),
  .ZN(_0083_)
);

INV_X1 _1808_ (
  .A(_1107_),
  .ZN(_0084_)
);

XNOR2_X1 _1809_ (
  .A(_0083_),
  .B(_0084_),
  .ZN(_0085_)
);

OAI21_X1 _1810_ (
  .A(_0076_),
  .B1(_0085_),
  .B2(_0581_),
  .ZN(_0086_)
);

NAND2_X1 _1811_ (
  .A1(_0387_),
  .A2(result[9]),
  .ZN(_0087_)
);

NAND2_X1 _1812_ (
  .A1(_0086_),
  .A2(_0087_),
  .ZN(_0028_)
);

NAND2_X1 _1813_ (
  .A1(_0385_),
  .A2(result[10]),
  .ZN(_0088_)
);

OAI21_X1 _1814_ (
  .A(_0632_),
  .B1(_0611_),
  .B2(_0634_),
  .ZN(_0089_)
);

NAND2_X1 _1815_ (
  .A1(_1105_),
  .A2(_1107_),
  .ZN(_0090_)
);

NOR2_X1 _1816_ (
  .A1(_0065_),
  .A2(_0090_),
  .ZN(_0091_)
);

NAND2_X1 _1817_ (
  .A1(_0089_),
  .A2(_0091_),
  .ZN(_0092_)
);

INV_X1 _1818_ (
  .A(_1106_),
  .ZN(_0093_)
);

OAI21_X1 _1819_ (
  .A(_0093_),
  .B1(_0084_),
  .B2(_0080_),
  .ZN(_0094_)
);

INV_X1 _1820_ (
  .A(_0094_),
  .ZN(_0095_)
);

OAI21_X1 _1821_ (
  .A(_0095_),
  .B1(_0064_),
  .B2(_0090_),
  .ZN(_0096_)
);

INV_X1 _1822_ (
  .A(_0096_),
  .ZN(_0097_)
);

NOR3_X1 _1823_ (
  .A1(_0634_),
  .A2(_0589_),
  .A3(_0609_),
  .ZN(_0098_)
);

INV_X1 _1824_ (
  .A(_0679_),
  .ZN(_0099_)
);

NAND3_X1 _1825_ (
  .A1(_0098_),
  .A2(_0099_),
  .A3(_0091_),
  .ZN(_0100_)
);

NAND3_X1 _1826_ (
  .A1(_0092_),
  .A2(_0097_),
  .A3(_0100_),
  .ZN(_0101_)
);

INV_X1 _1827_ (
  .A(_1109_),
  .ZN(_0102_)
);

XNOR2_X1 _1828_ (
  .A(_0101_),
  .B(_0102_),
  .ZN(_0103_)
);

NOR2_X1 _1829_ (
  .A1(_0103_),
  .A2(_0581_),
  .ZN(_0104_)
);

OAI21_X1 _1830_ (
  .A(_0368_),
  .B1(_0584_),
  .B2(\ext_mult_res[10] ),
  .ZN(_0105_)
);

OAI21_X1 _1831_ (
  .A(_0088_),
  .B1(_0104_),
  .B2(_0105_),
  .ZN(_0029_)
);

NAND2_X1 _1832_ (
  .A1(_0385_),
  .A2(result[11]),
  .ZN(_0106_)
);

NAND2_X1 _1833_ (
  .A1(_1107_),
  .A2(_1109_),
  .ZN(_0107_)
);

NOR2_X2 _1834_ (
  .A1(_0077_),
  .A2(_0107_),
  .ZN(_0108_)
);

NAND2_X1 _1835_ (
  .A1(_0051_),
  .A2(_0108_),
  .ZN(_0109_)
);

INV_X1 _1836_ (
  .A(_1108_),
  .ZN(_0110_)
);

OAI21_X1 _1837_ (
  .A(_0110_),
  .B1(_0102_),
  .B2(_0093_),
  .ZN(_0111_)
);

INV_X1 _1838_ (
  .A(_0111_),
  .ZN(_0112_)
);

OAI21_X1 _1839_ (
  .A(_0112_),
  .B1(_0082_),
  .B2(_0107_),
  .ZN(_0113_)
);

INV_X1 _1840_ (
  .A(_0113_),
  .ZN(_0114_)
);

NAND2_X1 _1841_ (
  .A1(_0109_),
  .A2(_0114_),
  .ZN(_0115_)
);

INV_X1 _1842_ (
  .A(_0115_),
  .ZN(_0116_)
);

NAND4_X1 _1843_ (
  .A1(_0108_),
  .A2(_0618_),
  .A3(_0636_),
  .A4(_0624_),
  .ZN(_0117_)
);

INV_X1 _1844_ (
  .A(_0117_),
  .ZN(_0118_)
);

INV_X1 _1845_ (
  .A(_0602_),
  .ZN(_0119_)
);

NAND2_X1 _1846_ (
  .A1(_0118_),
  .A2(_0119_),
  .ZN(_0120_)
);

NAND2_X1 _1847_ (
  .A1(_0116_),
  .A2(_0120_),
  .ZN(_0121_)
);

INV_X1 _1848_ (
  .A(_1111_),
  .ZN(_0122_)
);

NAND2_X1 _1849_ (
  .A1(_0121_),
  .A2(_0122_),
  .ZN(_0123_)
);

NAND3_X1 _1850_ (
  .A1(_0116_),
  .A2(_1111_),
  .A3(_0120_),
  .ZN(_0124_)
);

NAND3_X1 _1851_ (
  .A1(_0123_),
  .A2(_0124_),
  .A3(_0604_),
  .ZN(_0125_)
);

NAND2_X1 _1852_ (
  .A1(_0125_),
  .A2(_0374_),
  .ZN(_0126_)
);

NOR2_X1 _1853_ (
  .A1(_0584_),
  .A2(\ext_mult_res[11] ),
  .ZN(_0127_)
);

OAI21_X1 _1854_ (
  .A(_0106_),
  .B1(_0126_),
  .B2(_0127_),
  .ZN(_0030_)
);

NAND2_X1 _1855_ (
  .A1(_0385_),
  .A2(result[12]),
  .ZN(_0128_)
);

NAND2_X1 _1856_ (
  .A1(_1109_),
  .A2(_1111_),
  .ZN(_0129_)
);

NOR2_X1 _1857_ (
  .A1(_0090_),
  .A2(_0129_),
  .ZN(_0130_)
);

NAND2_X1 _1858_ (
  .A1(_0066_),
  .A2(_0130_),
  .ZN(_0131_)
);

INV_X1 _1859_ (
  .A(_1110_),
  .ZN(_0132_)
);

OAI21_X1 _1860_ (
  .A(_0132_),
  .B1(_0122_),
  .B2(_0110_),
  .ZN(_0133_)
);

INV_X1 _1861_ (
  .A(_0133_),
  .ZN(_0134_)
);

OAI21_X1 _1862_ (
  .A(_0134_),
  .B1(_0095_),
  .B2(_0129_),
  .ZN(_0135_)
);

INV_X1 _1863_ (
  .A(_0135_),
  .ZN(_0136_)
);

NAND2_X1 _1864_ (
  .A1(_0131_),
  .A2(_0136_),
  .ZN(_0137_)
);

INV_X1 _1865_ (
  .A(_0137_),
  .ZN(_0138_)
);

NAND2_X1 _1866_ (
  .A1(_0068_),
  .A2(_0130_),
  .ZN(_0139_)
);

INV_X1 _1867_ (
  .A(_0139_),
  .ZN(_0140_)
);

NAND2_X1 _1868_ (
  .A1(_0612_),
  .A2(_0140_),
  .ZN(_0141_)
);

NAND2_X1 _1869_ (
  .A1(_0138_),
  .A2(_0141_),
  .ZN(_0142_)
);

INV_X1 _1870_ (
  .A(_1113_),
  .ZN(_0143_)
);

NAND2_X1 _1871_ (
  .A1(_0142_),
  .A2(_0143_),
  .ZN(_0144_)
);

NAND3_X1 _1872_ (
  .A1(_0138_),
  .A2(_1113_),
  .A3(_0141_),
  .ZN(_0145_)
);

AND3_X1 _1873_ (
  .A1(_0144_),
  .A2(_0145_),
  .A3(_0594_),
  .ZN(_0146_)
);

OAI21_X1 _1874_ (
  .A(_0368_),
  .B1(_0584_),
  .B2(\ext_mult_res[12] ),
  .ZN(_0147_)
);

OAI21_X1 _1875_ (
  .A(_0128_),
  .B1(_0146_),
  .B2(_0147_),
  .ZN(_0031_)
);

NAND2_X1 _1876_ (
  .A1(_0385_),
  .A2(result[13]),
  .ZN(_0148_)
);

NAND2_X1 _1877_ (
  .A1(_0048_),
  .A2(_0078_),
  .ZN(_0149_)
);

NAND2_X1 _1878_ (
  .A1(_0082_),
  .A2(_0149_),
  .ZN(_0150_)
);

NAND2_X1 _1879_ (
  .A1(_1111_),
  .A2(_1113_),
  .ZN(_0151_)
);

NOR2_X1 _1880_ (
  .A1(_0107_),
  .A2(_0151_),
  .ZN(_0152_)
);

NAND2_X1 _1881_ (
  .A1(_0150_),
  .A2(_0152_),
  .ZN(_0153_)
);

INV_X1 _1882_ (
  .A(_0151_),
  .ZN(_0154_)
);

NAND2_X1 _1883_ (
  .A1(_0111_),
  .A2(_0154_),
  .ZN(_0155_)
);

INV_X1 _1884_ (
  .A(_1112_),
  .ZN(_0156_)
);

OAI21_X1 _1885_ (
  .A(_0156_),
  .B1(_0143_),
  .B2(_0132_),
  .ZN(_0157_)
);

INV_X1 _1886_ (
  .A(_0157_),
  .ZN(_0158_)
);

NAND2_X1 _1887_ (
  .A1(_0155_),
  .A2(_0158_),
  .ZN(_0159_)
);

INV_X1 _1888_ (
  .A(_0159_),
  .ZN(_0160_)
);

NAND2_X1 _1889_ (
  .A1(_0153_),
  .A2(_0160_),
  .ZN(_0161_)
);

INV_X1 _1890_ (
  .A(_0161_),
  .ZN(_0162_)
);

INV_X1 _1891_ (
  .A(_0623_),
  .ZN(_0163_)
);

NOR2_X2 _1892_ (
  .A1(_0050_),
  .A2(_0077_),
  .ZN(_0164_)
);

NAND2_X1 _1893_ (
  .A1(_0164_),
  .A2(_0152_),
  .ZN(_0165_)
);

OAI21_X1 _1894_ (
  .A(_0162_),
  .B1(_0163_),
  .B2(_0165_),
  .ZN(_0166_)
);

INV_X1 _1895_ (
  .A(_1115_),
  .ZN(_0167_)
);

XNOR2_X1 _1896_ (
  .A(_0166_),
  .B(_0167_),
  .ZN(_0168_)
);

NOR2_X1 _1897_ (
  .A1(_0168_),
  .A2(_0581_),
  .ZN(_0169_)
);

OAI21_X1 _1898_ (
  .A(_0368_),
  .B1(_0604_),
  .B2(\ext_mult_res[13] ),
  .ZN(_0170_)
);

OAI21_X1 _1899_ (
  .A(_0148_),
  .B1(_0169_),
  .B2(_0170_),
  .ZN(_0032_)
);

NAND2_X1 _1900_ (
  .A1(_1113_),
  .A2(_1115_),
  .ZN(_0171_)
);

NOR2_X1 _1901_ (
  .A1(_0129_),
  .A2(_0171_),
  .ZN(_0172_)
);

NAND3_X1 _1902_ (
  .A1(_0635_),
  .A2(_0091_),
  .A3(_0172_),
  .ZN(_0173_)
);

INV_X1 _1903_ (
  .A(_1114_),
  .ZN(_0174_)
);

OAI21_X1 _1904_ (
  .A(_0174_),
  .B1(_0167_),
  .B2(_0156_),
  .ZN(_0175_)
);

INV_X1 _1905_ (
  .A(_0175_),
  .ZN(_0176_)
);

OAI21_X1 _1906_ (
  .A(_0176_),
  .B1(_0134_),
  .B2(_0171_),
  .ZN(_0177_)
);

AOI21_X1 _1907_ (
  .A(_0177_),
  .B1(_0172_),
  .B2(_0096_),
  .ZN(_0178_)
);

NAND2_X1 _1908_ (
  .A1(_0173_),
  .A2(_0178_),
  .ZN(_0179_)
);

INV_X1 _1909_ (
  .A(_1117_),
  .ZN(_0180_)
);

NAND2_X1 _1910_ (
  .A1(_0179_),
  .A2(_0180_),
  .ZN(_0181_)
);

NAND3_X1 _1911_ (
  .A1(_0173_),
  .A2(_1117_),
  .A3(_0178_),
  .ZN(_0182_)
);

NAND3_X1 _1912_ (
  .A1(_0181_),
  .A2(_0182_),
  .A3(_0604_),
  .ZN(_0183_)
);

OAI21_X1 _1913_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[14] ),
  .ZN(_0184_)
);

INV_X1 _1914_ (
  .A(_0184_),
  .ZN(_0185_)
);

NAND2_X1 _1915_ (
  .A1(_0183_),
  .A2(_0185_),
  .ZN(_0186_)
);

NAND2_X1 _1916_ (
  .A1(_0387_),
  .A2(result[14]),
  .ZN(_0187_)
);

NAND2_X1 _1917_ (
  .A1(_0186_),
  .A2(_0187_),
  .ZN(_0033_)
);

NAND2_X1 _1918_ (
  .A1(_1115_),
  .A2(_1117_),
  .ZN(_0188_)
);

NOR2_X1 _1919_ (
  .A1(_0151_),
  .A2(_0188_),
  .ZN(_0189_)
);

NAND3_X1 _1920_ (
  .A1(_0053_),
  .A2(_0108_),
  .A3(_0189_),
  .ZN(_0190_)
);

INV_X1 _1921_ (
  .A(_1116_),
  .ZN(_0191_)
);

OAI21_X1 _1922_ (
  .A(_0191_),
  .B1(_0180_),
  .B2(_0174_),
  .ZN(_0192_)
);

INV_X1 _1923_ (
  .A(_0192_),
  .ZN(_0193_)
);

OAI21_X1 _1924_ (
  .A(_0193_),
  .B1(_0158_),
  .B2(_0188_),
  .ZN(_0194_)
);

AOI21_X1 _1925_ (
  .A(_0194_),
  .B1(_0189_),
  .B2(_0113_),
  .ZN(_0195_)
);

NAND2_X1 _1926_ (
  .A1(_0190_),
  .A2(_0195_),
  .ZN(_0196_)
);

INV_X1 _1927_ (
  .A(_1119_),
  .ZN(_0197_)
);

NAND2_X1 _1928_ (
  .A1(_0196_),
  .A2(_0197_),
  .ZN(_0198_)
);

NAND3_X1 _1929_ (
  .A1(_0190_),
  .A2(_1119_),
  .A3(_0195_),
  .ZN(_0199_)
);

NAND3_X1 _1930_ (
  .A1(_0198_),
  .A2(_0199_),
  .A3(_0604_),
  .ZN(_0200_)
);

OAI21_X1 _1931_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[15] ),
  .ZN(_0201_)
);

INV_X1 _1932_ (
  .A(_0201_),
  .ZN(_0202_)
);

NAND2_X1 _1933_ (
  .A1(_0200_),
  .A2(_0202_),
  .ZN(_0203_)
);

NAND2_X1 _1934_ (
  .A1(_0387_),
  .A2(result[15]),
  .ZN(_0204_)
);

NAND2_X1 _1935_ (
  .A1(_0203_),
  .A2(_0204_),
  .ZN(_0034_)
);

OAI21_X1 _1936_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[16] ),
  .ZN(_0205_)
);

INV_X1 _1937_ (
  .A(_0205_),
  .ZN(_0206_)
);

NAND2_X1 _1938_ (
  .A1(_1117_),
  .A2(_1119_),
  .ZN(_0207_)
);

NOR2_X1 _1939_ (
  .A1(_0171_),
  .A2(_0207_),
  .ZN(_0208_)
);

NAND3_X1 _1940_ (
  .A1(_0070_),
  .A2(_0130_),
  .A3(_0208_),
  .ZN(_0209_)
);

BUF_X2 _1941_ (
  .A(_1121_),
  .Z(_0210_)
);

INV_X1 _1942_ (
  .A(_1118_),
  .ZN(_0211_)
);

OAI21_X1 _1943_ (
  .A(_0211_),
  .B1(_0197_),
  .B2(_0191_),
  .ZN(_0212_)
);

INV_X1 _1944_ (
  .A(_0212_),
  .ZN(_0213_)
);

OAI21_X1 _1945_ (
  .A(_0213_),
  .B1(_0176_),
  .B2(_0207_),
  .ZN(_0214_)
);

AOI21_X1 _1946_ (
  .A(_0214_),
  .B1(_0208_),
  .B2(_0135_),
  .ZN(_0215_)
);

NAND3_X1 _1947_ (
  .A1(_0209_),
  .A2(_0210_),
  .A3(_0215_),
  .ZN(_0216_)
);

NAND2_X1 _1948_ (
  .A1(_0216_),
  .A2(_0604_),
  .ZN(_0217_)
);

AOI21_X1 _1949_ (
  .A(_0210_),
  .B1(_0209_),
  .B2(_0215_),
  .ZN(_0218_)
);

OAI21_X1 _1950_ (
  .A(_0206_),
  .B1(_0217_),
  .B2(_0218_),
  .ZN(_0219_)
);

NAND2_X1 _1951_ (
  .A1(_0387_),
  .A2(result[16]),
  .ZN(_0220_)
);

NAND2_X1 _1952_ (
  .A1(_0219_),
  .A2(_0220_),
  .ZN(_0035_)
);

OAI21_X1 _1953_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[17] ),
  .ZN(_0221_)
);

INV_X1 _1954_ (
  .A(_0221_),
  .ZN(_0222_)
);

OAI21_X1 _1955_ (
  .A(_0599_),
  .B1(_0589_),
  .B2(_0598_),
  .ZN(_0223_)
);

INV_X1 _1956_ (
  .A(_0223_),
  .ZN(_0224_)
);

OAI21_X1 _1957_ (
  .A(_0622_),
  .B1(_0224_),
  .B2(_0617_),
  .ZN(_0225_)
);

NAND2_X1 _1958_ (
  .A1(_0225_),
  .A2(_0164_),
  .ZN(_0226_)
);

INV_X1 _1959_ (
  .A(_0150_),
  .ZN(_0227_)
);

NAND2_X1 _1960_ (
  .A1(_0226_),
  .A2(_0227_),
  .ZN(_0228_)
);

NAND2_X2 _1961_ (
  .A1(_1119_),
  .A2(_0210_),
  .ZN(_0229_)
);

NOR2_X2 _1962_ (
  .A1(_0188_),
  .A2(_0229_),
  .ZN(_0230_)
);

AND2_X1 _1963_ (
  .A1(_0152_),
  .A2(_0230_),
  .ZN(_0231_)
);

NAND2_X1 _1964_ (
  .A1(_0228_),
  .A2(_0231_),
  .ZN(_0232_)
);

INV_X1 _1965_ (
  .A(_0229_),
  .ZN(_0233_)
);

NAND2_X1 _1966_ (
  .A1(_0192_),
  .A2(_0233_),
  .ZN(_0234_)
);

INV_X1 _1967_ (
  .A(_1120_),
  .ZN(_0235_)
);

INV_X1 _1968_ (
  .A(_0210_),
  .ZN(_0236_)
);

OAI21_X1 _1969_ (
  .A(_0235_),
  .B1(_0236_),
  .B2(_0211_),
  .ZN(_0237_)
);

INV_X1 _1970_ (
  .A(_0237_),
  .ZN(_0238_)
);

NAND2_X1 _1971_ (
  .A1(_0234_),
  .A2(_0238_),
  .ZN(_0239_)
);

AOI21_X1 _1972_ (
  .A(_0239_),
  .B1(_0230_),
  .B2(_0159_),
  .ZN(_0240_)
);

AND3_X1 _1973_ (
  .A1(_0618_),
  .A2(_1091_),
  .A3(_1093_),
  .ZN(_0241_)
);

NAND4_X1 _1974_ (
  .A1(_0231_),
  .A2(_0241_),
  .A3(_0164_),
  .A4(_1088_),
  .ZN(_0242_)
);

NAND3_X1 _1975_ (
  .A1(_0232_),
  .A2(_0240_),
  .A3(_0242_),
  .ZN(_0243_)
);

INV_X1 _1976_ (
  .A(_1123_),
  .ZN(_0244_)
);

NAND2_X1 _1977_ (
  .A1(_0243_),
  .A2(_0244_),
  .ZN(_0245_)
);

NAND2_X1 _1978_ (
  .A1(_0245_),
  .A2(_0604_),
  .ZN(_0246_)
);

NOR2_X1 _1979_ (
  .A1(_0243_),
  .A2(_0244_),
  .ZN(_0247_)
);

OAI21_X1 _1980_ (
  .A(_0222_),
  .B1(_0246_),
  .B2(_0247_),
  .ZN(_0248_)
);

NAND2_X1 _1981_ (
  .A1(_0387_),
  .A2(result[17]),
  .ZN(_0249_)
);

NAND2_X1 _1982_ (
  .A1(_0248_),
  .A2(_0249_),
  .ZN(_0036_)
);

NOR2_X1 _1983_ (
  .A1(_0368_),
  .A2(result[18]),
  .ZN(_0250_)
);

NAND2_X1 _1984_ (
  .A1(_0092_),
  .A2(_0097_),
  .ZN(_0251_)
);

NAND2_X1 _1985_ (
  .A1(_0210_),
  .A2(_1123_),
  .ZN(_0252_)
);

NOR2_X1 _1986_ (
  .A1(_0207_),
  .A2(_0252_),
  .ZN(_0253_)
);

AND2_X1 _1987_ (
  .A1(_0172_),
  .A2(_0253_),
  .ZN(_0254_)
);

NAND2_X1 _1988_ (
  .A1(_0251_),
  .A2(_0254_),
  .ZN(_0255_)
);

INV_X1 _1989_ (
  .A(_1122_),
  .ZN(_0256_)
);

OAI21_X1 _1990_ (
  .A(_0256_),
  .B1(_0244_),
  .B2(_0235_),
  .ZN(_0257_)
);

INV_X1 _1991_ (
  .A(_0257_),
  .ZN(_0258_)
);

OAI21_X1 _1992_ (
  .A(_0258_),
  .B1(_0213_),
  .B2(_0252_),
  .ZN(_0259_)
);

AOI21_X1 _1993_ (
  .A(_0259_),
  .B1(_0253_),
  .B2(_0177_),
  .ZN(_0260_)
);

NAND4_X1 _1994_ (
  .A1(_0254_),
  .A2(_0091_),
  .A3(_0098_),
  .A4(_0099_),
  .ZN(_0261_)
);

NAND3_X1 _1995_ (
  .A1(_0255_),
  .A2(_0260_),
  .A3(_0261_),
  .ZN(_0262_)
);

NAND2_X1 _1996_ (
  .A1(_0262_),
  .A2(_1125_),
  .ZN(_0263_)
);

INV_X1 _1997_ (
  .A(_1125_),
  .ZN(_0264_)
);

NAND4_X1 _1998_ (
  .A1(_0255_),
  .A2(_0260_),
  .A3(_0264_),
  .A4(_0261_),
  .ZN(_0265_)
);

NAND3_X1 _1999_ (
  .A1(_0263_),
  .A2(_0265_),
  .A3(_0584_),
  .ZN(_0266_)
);

NAND2_X1 _2000_ (
  .A1(_0581_),
  .A2(\ext_mult_res[18] ),
  .ZN(_0267_)
);

NAND2_X1 _2001_ (
  .A1(_0267_),
  .A2(_0371_),
  .ZN(_0268_)
);

INV_X1 _2002_ (
  .A(_0268_),
  .ZN(_0269_)
);

AOI21_X1 _2003_ (
  .A(_0250_),
  .B1(_0266_),
  .B2(_0269_),
  .ZN(_0037_)
);

NOR2_X1 _2004_ (
  .A1(_0368_),
  .A2(result[19]),
  .ZN(_0270_)
);

NAND2_X1 _2005_ (
  .A1(_1123_),
  .A2(_1125_),
  .ZN(_0271_)
);

NOR2_X1 _2006_ (
  .A1(_0229_),
  .A2(_0271_),
  .ZN(_0272_)
);

AND2_X1 _2007_ (
  .A1(_0189_),
  .A2(_0272_),
  .ZN(_0273_)
);

NAND2_X1 _2008_ (
  .A1(_0115_),
  .A2(_0273_),
  .ZN(_0274_)
);

INV_X1 _2009_ (
  .A(_1124_),
  .ZN(_0275_)
);

OAI21_X1 _2010_ (
  .A(_0275_),
  .B1(_0264_),
  .B2(_0256_),
  .ZN(_0276_)
);

INV_X1 _2011_ (
  .A(_0276_),
  .ZN(_0277_)
);

OAI21_X1 _2012_ (
  .A(_0277_),
  .B1(_0238_),
  .B2(_0271_),
  .ZN(_0278_)
);

AOI21_X1 _2013_ (
  .A(_0278_),
  .B1(_0272_),
  .B2(_0194_),
  .ZN(_0279_)
);

NAND3_X1 _2014_ (
  .A1(_0118_),
  .A2(_0119_),
  .A3(_0273_),
  .ZN(_0280_)
);

NAND3_X1 _2015_ (
  .A1(_0274_),
  .A2(_0279_),
  .A3(_0280_),
  .ZN(_0281_)
);

NAND2_X1 _2016_ (
  .A1(_0281_),
  .A2(_1127_),
  .ZN(_0282_)
);

INV_X1 _2017_ (
  .A(_1127_),
  .ZN(_0283_)
);

NAND4_X1 _2018_ (
  .A1(_0274_),
  .A2(_0279_),
  .A3(_0283_),
  .A4(_0280_),
  .ZN(_0284_)
);

NAND3_X1 _2019_ (
  .A1(_0282_),
  .A2(_0284_),
  .A3(_0584_),
  .ZN(_0285_)
);

AOI21_X1 _2020_ (
  .A(_0270_),
  .B1(_0285_),
  .B2(_0269_),
  .ZN(_0038_)
);

NOR2_X1 _2021_ (
  .A1(_0368_),
  .A2(result[20]),
  .ZN(_0286_)
);

NAND2_X1 _2022_ (
  .A1(_1125_),
  .A2(_1127_),
  .ZN(_0287_)
);

NOR2_X1 _2023_ (
  .A1(_0252_),
  .A2(_0287_),
  .ZN(_0288_)
);

AND2_X1 _2024_ (
  .A1(_0208_),
  .A2(_0288_),
  .ZN(_0289_)
);

NAND2_X1 _2025_ (
  .A1(_0137_),
  .A2(_0289_),
  .ZN(_0290_)
);

INV_X1 _2026_ (
  .A(_1126_),
  .ZN(_0291_)
);

OAI21_X1 _2027_ (
  .A(_0291_),
  .B1(_0283_),
  .B2(_0275_),
  .ZN(_0292_)
);

INV_X1 _2028_ (
  .A(_0292_),
  .ZN(_0293_)
);

OAI21_X1 _2029_ (
  .A(_0293_),
  .B1(_0258_),
  .B2(_0287_),
  .ZN(_0294_)
);

AOI21_X1 _2030_ (
  .A(_0294_),
  .B1(_0288_),
  .B2(_0214_),
  .ZN(_0295_)
);

NAND3_X1 _2031_ (
  .A1(_0612_),
  .A2(_0140_),
  .A3(_0289_),
  .ZN(_0296_)
);

NAND3_X1 _2032_ (
  .A1(_0290_),
  .A2(_0295_),
  .A3(_0296_),
  .ZN(_0297_)
);

NAND2_X1 _2033_ (
  .A1(_0297_),
  .A2(_1129_),
  .ZN(_0298_)
);

INV_X1 _2034_ (
  .A(_1129_),
  .ZN(_0299_)
);

NAND4_X1 _2035_ (
  .A1(_0290_),
  .A2(_0295_),
  .A3(_0299_),
  .A4(_0296_),
  .ZN(_0300_)
);

NAND3_X1 _2036_ (
  .A1(_0298_),
  .A2(_0300_),
  .A3(_0584_),
  .ZN(_0301_)
);

AOI21_X1 _2037_ (
  .A(_0286_),
  .B1(_0301_),
  .B2(_0269_),
  .ZN(_0039_)
);

NAND2_X1 _2038_ (
  .A1(_1127_),
  .A2(_1129_),
  .ZN(_0302_)
);

NOR2_X1 _2039_ (
  .A1(_0271_),
  .A2(_0302_),
  .ZN(_0303_)
);

NAND2_X1 _2040_ (
  .A1(_0230_),
  .A2(_0303_),
  .ZN(_0304_)
);

INV_X1 _2041_ (
  .A(_0304_),
  .ZN(_0305_)
);

NAND2_X1 _2042_ (
  .A1(_0161_),
  .A2(_0305_),
  .ZN(_0306_)
);

INV_X1 _2043_ (
  .A(_0303_),
  .ZN(_0307_)
);

AOI21_X1 _2044_ (
  .A(_0307_),
  .B1(_0234_),
  .B2(_0238_),
  .ZN(_0308_)
);

INV_X1 _2045_ (
  .A(_1128_),
  .ZN(_0309_)
);

OAI21_X1 _2046_ (
  .A(_0309_),
  .B1(_0299_),
  .B2(_0291_),
  .ZN(_0310_)
);

INV_X1 _2047_ (
  .A(_0310_),
  .ZN(_0311_)
);

OAI21_X1 _2048_ (
  .A(_0311_),
  .B1(_0277_),
  .B2(_0302_),
  .ZN(_0312_)
);

NOR2_X1 _2049_ (
  .A1(_0308_),
  .A2(_0312_),
  .ZN(_0313_)
);

NOR2_X1 _2050_ (
  .A1(_0165_),
  .A2(_0304_),
  .ZN(_0314_)
);

NAND2_X1 _2051_ (
  .A1(_0623_),
  .A2(_0314_),
  .ZN(_0315_)
);

XOR2_X1 _2052_ (
  .A(\ext_mult_res[18] ),
  .B(result[21]),
  .Z(_0316_)
);

NAND4_X1 _2053_ (
  .A1(_0306_),
  .A2(_0313_),
  .A3(_0315_),
  .A4(_0316_),
  .ZN(_0317_)
);

NAND3_X1 _2054_ (
  .A1(_0306_),
  .A2(_0313_),
  .A3(_0315_),
  .ZN(_0318_)
);

INV_X1 _2055_ (
  .A(_0316_),
  .ZN(_0319_)
);

NAND2_X1 _2056_ (
  .A1(_0318_),
  .A2(_0319_),
  .ZN(_0320_)
);

NAND2_X1 _2057_ (
  .A1(_0317_),
  .A2(_0320_),
  .ZN(_0321_)
);

NAND2_X1 _2058_ (
  .A1(_0321_),
  .A2(_0594_),
  .ZN(_0322_)
);

NAND2_X1 _2059_ (
  .A1(_0322_),
  .A2(_0267_),
  .ZN(_0323_)
);

NAND2_X1 _2060_ (
  .A1(_0323_),
  .A2(_0372_),
  .ZN(_0324_)
);

NAND2_X1 _2061_ (
  .A1(_0387_),
  .A2(result[21]),
  .ZN(_0325_)
);

NAND2_X1 _2062_ (
  .A1(_0324_),
  .A2(_0325_),
  .ZN(_0040_)
);

FA_X1 _2063_ (
  .A(_0676_),
  .B(_0677_),
  .CI(_0678_),
  .CO(_0679_),
  .S(_0680_)
);

FA_X1 _2064_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0684_),
  .S(_0685_)
);

FA_X1 _2065_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0689_),
  .S(_0690_)
);

FA_X1 _2066_ (
  .A(_0690_),
  .B(_0684_),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0692_),
  .S(_0693_)
);

FA_X1 _2067_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0697_),
  .S(_0698_)
);

FA_X1 _2068_ (
  .A(_0698_),
  .B(_0699_),
  .CI(_0700_),
  .CO(_0701_),
  .S(_0702_)
);

FA_X1 _2069_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0706_),
  .S(_0707_)
);

FA_X1 _2070_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0711_),
  .S(_0712_)
);

FA_X1 _2071_ (
  .A(_0707_),
  .B(_0697_),
  .CI(_0712_),
  .CO(_0713_),
  .S(_0714_)
);

FA_X1 _2072_ (
  .A(_0715_),
  .B(_0716_),
  .CI(_0717_),
  .CO(_0718_),
  .S(_0719_)
);

FA_X1 _2073_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0723_),
  .S(_0724_)
);

FA_X1 _2074_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0728_),
  .S(_0729_)
);

FA_X1 _2075_ (
  .A(_0724_),
  .B(_0706_),
  .CI(_0729_),
  .CO(_0730_),
  .S(_0731_)
);

FA_X1 _2076_ (
  .A(_0731_),
  .B(_0713_),
  .CI(_0732_),
  .CO(_0733_),
  .S(_0734_)
);

FA_X1 _2077_ (
  .A(_0735_),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0738_),
  .S(_0739_)
);

FA_X1 _2078_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0743_),
  .S(_0744_)
);

FA_X1 _2079_ (
  .A(_0744_),
  .B(_0739_),
  .CI(_0745_),
  .CO(_0746_),
  .S(_0747_)
);

FA_X1 _2080_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0751_),
  .S(_0752_)
);

FA_X1 _2081_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0756_),
  .S(_0757_)
);

FA_X1 _2082_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0761_),
  .S(_0762_)
);

FA_X1 _2083_ (
  .A(_0765_),
  .B(_0766_),
  .CI(_0767_),
  .CO(_0768_),
  .S(_0769_)
);

FA_X1 _2084_ (
  .A(_0770_),
  .B(_0747_),
  .CI(_0771_),
  .CO(_0772_),
  .S(_0773_)
);

FA_X1 _2085_ (
  .A(_0757_),
  .B(_0774_),
  .CI(_0775_),
  .CO(_0776_),
  .S(_0777_)
);

FA_X1 _2086_ (
  .A(_0778_),
  .B(_0779_),
  .CI(_0780_),
  .CO(_0781_),
  .S(_0782_)
);

FA_X1 _2087_ (
  .A(_0777_),
  .B(_0730_),
  .CI(_0784_),
  .CO(_0783_),
  .S(_0785_)
);

FA_X1 _2088_ (
  .A(_0786_),
  .B(_0733_),
  .CI(_0787_),
  .CO(_0788_),
  .S(_0789_)
);

FA_X1 _2089_ (
  .A(_0790_),
  .B(_0791_),
  .CI(_0792_),
  .CO(_0793_),
  .S(_0794_)
);

FA_X1 _2090_ (
  .A(_0795_),
  .B(_0796_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0798_),
  .S(_0799_)
);

FA_X1 _2091_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0803_),
  .S(_0804_)
);

FA_X1 _2092_ (
  .A(_0799_),
  .B(_0738_),
  .CI(_0804_),
  .CO(_0805_),
  .S(_0806_)
);

FA_X1 _2093_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0809_),
  .S(_0810_)
);

FA_X1 _2094_ (
  .A(_0811_),
  .B(_0812_),
  .CI(_0813_),
  .CO(_0814_),
  .S(_0815_)
);

FA_X1 _2095_ (
  .A(_0806_),
  .B(_0746_),
  .CI(_0815_),
  .CO(_0816_),
  .S(_0817_)
);

FA_X1 _2096_ (
  .A(_0817_),
  .B(_0772_),
  .CI(_0818_),
  .CO(_0819_),
  .S(_0820_)
);

FA_X1 _2097_ (
  .A(_0821_),
  .B(_0822_),
  .CI(_0823_),
  .CO(_0824_),
  .S(_0825_)
);

FA_X1 _2098_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0829_),
  .S(_0830_)
);

FA_X1 _2099_ (
  .A(_0825_),
  .B(_0798_),
  .CI(_0830_),
  .CO(_0831_),
  .S(_0832_)
);

FA_X1 _2100_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0835_),
  .S(_0836_)
);

FA_X1 _2101_ (
  .A(_0837_),
  .B(_0838_),
  .CI(_0839_),
  .CO(_0840_),
  .S(_0841_)
);

FA_X1 _2102_ (
  .A(_0841_),
  .B(_0832_),
  .CI(_0805_),
  .CO(_0842_),
  .S(_0843_)
);

FA_X1 _2103_ (
  .A(_0816_),
  .B(_0843_),
  .CI(_0844_),
  .CO(_0845_),
  .S(_0846_)
);

FA_X1 _2104_ (
  .A(_0847_),
  .B(_0848_),
  .CI(_0849_),
  .CO(_0850_),
  .S(_0851_)
);

FA_X1 _2105_ (
  .A(_0852_),
  .B(_0853_),
  .CI(_0854_),
  .CO(_0855_),
  .S(_0856_)
);

FA_X1 _2106_ (
  .A(_0857_),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0860_),
  .S(_0861_)
);

FA_X1 _2107_ (
  .A(_0862_),
  .B(_0824_),
  .CI(_0861_),
  .CO(_0863_),
  .S(_0864_)
);

FA_X1 _2108_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0867_),
  .S(_0868_)
);

FA_X1 _2109_ (
  .A(_0829_),
  .B(_0868_),
  .CI(_0835_),
  .CO(_0869_),
  .S(_0870_)
);

FA_X1 _2110_ (
  .A(_0864_),
  .B(_0831_),
  .CI(_0870_),
  .CO(_0871_),
  .S(_0872_)
);

FA_X1 _2111_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0874_),
  .S(_0875_)
);

FA_X1 _2112_ (
  .A(_0872_),
  .B(_0842_),
  .CI(_0876_),
  .CO(_0877_),
  .S(_0878_)
);

FA_X1 _2113_ (
  .A(_0878_),
  .B(_0845_),
  .CI(_0879_),
  .CO(_0880_),
  .S(_0881_)
);

FA_X1 _2114_ (
  .A(_0852_),
  .B(_0882_),
  .CI(_0854_),
  .CO(_0883_),
  .S(_0884_)
);

FA_X1 _2115_ (
  .A(_0885_),
  .B(_0886_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0888_),
  .S(_0889_)
);

FA_X1 _2116_ (
  .A(_0890_),
  .B(_0891_),
  .CI(_0889_),
  .CO(_0892_),
  .S(_0893_)
);

FA_X1 _2117_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0896_),
  .S(_0897_)
);

FA_X1 _2118_ (
  .A(_0860_),
  .B(_0897_),
  .CI(_0867_),
  .CO(_0898_),
  .S(_0899_)
);

FA_X1 _2119_ (
  .A(_0893_),
  .B(_0863_),
  .CI(_0899_),
  .CO(_0900_),
  .S(_0901_)
);

FA_X1 _2120_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0902_),
  .S(_0903_)
);

FA_X1 _2121_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(_0904_),
  .CI(_0905_),
  .CO(_0906_),
  .S(_0907_)
);

FA_X1 _2122_ (
  .A(_0908_),
  .B(_0909_),
  .CI(_0910_),
  .CO(_0911_),
  .S(_0912_)
);

FA_X1 _2123_ (
  .A(_0901_),
  .B(_0871_),
  .CI(_0913_),
  .CO(_0914_),
  .S(_0915_)
);

FA_X1 _2124_ (
  .A(_0915_),
  .B(_0877_),
  .CI(_0916_),
  .CO(_0917_),
  .S(_0918_)
);

FA_X1 _2125_ (
  .A(_0919_),
  .B(_0920_),
  .CI(_0921_),
  .CO(_0922_),
  .S(_0923_)
);

FA_X1 _2126_ (
  .A(_0924_),
  .B(_0923_),
  .CI(_0890_),
  .CO(_0925_),
  .S(_0926_)
);

FA_X1 _2127_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0929_),
  .S(_0930_)
);

FA_X1 _2128_ (
  .A(_0888_),
  .B(_0930_),
  .CI(_0896_),
  .CO(_0931_),
  .S(_0932_)
);

FA_X1 _2129_ (
  .A(_0926_),
  .B(_0892_),
  .CI(_0932_),
  .CO(_0933_),
  .S(_0934_)
);

FA_X1 _2130_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0935_),
  .S(_0936_)
);

FA_X1 _2131_ (
  .A(_0937_),
  .B(_0938_),
  .CI(_0902_),
  .CO(_0939_),
  .S(_0940_)
);

FA_X1 _2132_ (
  .A(_0898_),
  .B(_0940_),
  .CI(_0906_),
  .CO(_0943_),
  .S(_0944_)
);

FA_X1 _2133_ (
  .A(_0934_),
  .B(_0900_),
  .CI(_0944_),
  .CO(_0945_),
  .S(_0946_)
);

FA_X1 _2134_ (
  .A(_0947_),
  .B(_0948_),
  .CI(_0911_),
  .CO(_0949_),
  .S(_0950_)
);

FA_X1 _2135_ (
  .A(_0951_),
  .B(_0952_),
  .CI(_0953_),
  .CO(_0954_),
  .S(_0955_)
);

FA_X1 _2136_ (
  .A(_0924_),
  .B(_0956_),
  .CI(_0890_),
  .CO(_0957_),
  .S(_0958_)
);

FA_X1 _2137_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(_0959_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0961_),
  .S(_0962_)
);

FA_X1 _2138_ (
  .A(_0922_),
  .B(_0962_),
  .CI(_0929_),
  .CO(_0963_),
  .S(_0964_)
);

FA_X1 _2139_ (
  .A(_0958_),
  .B(_0925_),
  .CI(_0964_),
  .CO(_0965_),
  .S(_0966_)
);

FA_X1 _2140_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0967_),
  .S(_0968_)
);

FA_X1 _2141_ (
  .A(_0969_),
  .B(_0970_),
  .CI(_0935_),
  .CO(_0971_),
  .S(_0972_)
);

FA_X1 _2142_ (
  .A(_0974_),
  .B(_0975_),
  .CI(_0976_),
  .CO(_0977_),
  .S(_0978_)
);

FA_X1 _2143_ (
  .A(_0966_),
  .B(_0933_),
  .CI(_0978_),
  .CO(_0979_),
  .S(_0980_)
);

FA_X1 _2144_ (
  .A(_0981_),
  .B(_0982_),
  .CI(_0983_),
  .CO(_0984_),
  .S(_0985_)
);

FA_X1 _2145_ (
  .A(_0951_),
  .B(_0986_),
  .CI(_0952_),
  .CO(_0987_),
  .S(_0988_)
);

FA_X1 _2146_ (
  .A(_0924_),
  .B(_0989_),
  .CI(_0890_),
  .CO(_0990_),
  .S(_0991_)
);

FA_X1 _2147_ (
  .A(_0992_),
  .B(_0993_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0994_),
  .S(_0995_)
);

FA_X1 _2148_ (
  .A(_0995_),
  .B(_0961_),
  .CI(_0996_),
  .CO(_0997_),
  .S(_0998_)
);

FA_X1 _2149_ (
  .A(_0998_),
  .B(_0991_),
  .CI(_0957_),
  .CO(_0999_),
  .S(_1000_)
);

FA_X1 _2150_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_1004_),
  .S(_1005_)
);

FA_X1 _2151_ (
  .A(_1005_),
  .B(_1006_),
  .CI(_0903_),
  .CO(_1007_),
  .S(_1008_)
);

FA_X1 _2152_ (
  .A(_1009_),
  .B(_1008_),
  .CI(_1010_),
  .CO(_1011_),
  .S(_1012_)
);

FA_X1 _2153_ (
  .A(_1000_),
  .B(_0965_),
  .CI(_1012_),
  .CO(_1013_),
  .S(_1014_)
);

FA_X1 _2154_ (
  .A(_1014_),
  .B(_0979_),
  .CI(_1015_),
  .CO(_1016_),
  .S(_1017_)
);

FA_X1 _2155_ (
  .A(_1018_),
  .B(_0984_),
  .CI(_1019_),
  .CO(_1020_),
  .S(_1021_)
);

FA_X1 _2156_ (
  .A(_1022_),
  .B(_1023_),
  .CI(_1024_),
  .CO(_1025_),
  .S(_1026_)
);

FA_X1 _2157_ (
  .A(_1027_),
  .B(_1028_),
  .CI(_0994_),
  .CO(_1029_),
  .S(_1030_)
);

FA_X1 _2158_ (
  .A(_0990_),
  .B(_1030_),
  .CI(_0991_),
  .CO(_1031_),
  .S(_1032_)
);

FA_X1 _2159_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_1034_),
  .S(_1035_)
);

FA_X1 _2160_ (
  .A(_1035_),
  .B(_1004_),
  .CI(_0936_),
  .CO(_1036_),
  .S(_1037_)
);

FA_X1 _2161_ (
  .A(_0997_),
  .B(_1038_),
  .CI(_1039_),
  .CO(_1040_),
  .S(_1041_)
);

FA_X1 _2162_ (
  .A(_1032_),
  .B(_0999_),
  .CI(_1041_),
  .CO(_1042_),
  .S(_1043_)
);

FA_X1 _2163_ (
  .A(_1043_),
  .B(_1013_),
  .CI(_1044_),
  .CO(_1045_),
  .S(_1046_)
);

FA_X1 _2164_ (
  .A(_1047_),
  .B(_1048_),
  .CI(_1049_),
  .CO(_1050_),
  .S(_1051_)
);

FA_X1 _2165_ (
  .A(_1052_),
  .B(_1053_),
  .CI(_1054_),
  .CO(_1055_),
  .S(_1056_)
);

FA_X1 _2166_ (
  .A(_1027_),
  .B(_1057_),
  .CI(_1058_),
  .CO(_1059_),
  .S(_1060_)
);

FA_X1 _2167_ (
  .A(_0990_),
  .B(_1060_),
  .CI(_0991_),
  .CO(_1061_),
  .S(_1062_)
);

FA_X1 _2168_ (
  .A(_0993_),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_1063_),
  .S(_1064_)
);

FA_X1 _2169_ (
  .A(_1034_),
  .B(_1064_),
  .CI(_0968_),
  .CO(_1065_),
  .S(_1066_)
);

FA_X1 _2170_ (
  .A(_1066_),
  .B(_1036_),
  .CI(_1067_),
  .CO(_1068_),
  .S(_1069_)
);

FA_X1 _2171_ (
  .A(_1069_),
  .B(_1062_),
  .CI(_1031_),
  .CO(_1070_),
  .S(_1071_)
);

FA_X1 _2172_ (
  .A(_0973_),
  .B(_0875_),
  .CI(_1072_),
  .CO(_1073_),
  .S(_1074_)
);

FA_X1 _2173_ (
  .A(_1075_),
  .B(_1076_),
  .CI(_1077_),
  .CO(_1078_),
  .S(_1079_)
);

FA_X1 _2174_ (
  .A(_1071_),
  .B(_1042_),
  .CI(_1080_),
  .CO(_1081_),
  .S(_1082_)
);

FA_X1 _2175_ (
  .A(_1083_),
  .B(_1084_),
  .CI(_1085_),
  .CO(_1086_),
  .S(_1087_)
);

HA_X1 _2176_ (
  .A(result[0]),
  .B(\ext_mult_res[0] ),
  .CO(_1088_),
  .S(_1089_)
);

HA_X1 _2177_ (
  .A(result[1]),
  .B(\ext_mult_res[1] ),
  .CO(_1090_),
  .S(_1091_)
);

HA_X1 _2178_ (
  .A(result[2]),
  .B(\ext_mult_res[2] ),
  .CO(_1092_),
  .S(_1093_)
);

HA_X1 _2179_ (
  .A(result[3]),
  .B(\ext_mult_res[3] ),
  .CO(_1094_),
  .S(_1095_)
);

HA_X1 _2180_ (
  .A(result[4]),
  .B(\ext_mult_res[4] ),
  .CO(_1096_),
  .S(_1097_)
);

HA_X1 _2181_ (
  .A(result[5]),
  .B(\ext_mult_res[5] ),
  .CO(_1098_),
  .S(_1099_)
);

HA_X1 _2182_ (
  .A(result[6]),
  .B(\ext_mult_res[6] ),
  .CO(_1100_),
  .S(_1101_)
);

HA_X1 _2183_ (
  .A(result[7]),
  .B(\ext_mult_res[7] ),
  .CO(_1102_),
  .S(_1103_)
);

HA_X1 _2184_ (
  .A(result[8]),
  .B(\ext_mult_res[8] ),
  .CO(_1104_),
  .S(_1105_)
);

HA_X1 _2185_ (
  .A(result[9]),
  .B(\ext_mult_res[9] ),
  .CO(_1106_),
  .S(_1107_)
);

HA_X1 _2186_ (
  .A(result[10]),
  .B(\ext_mult_res[10] ),
  .CO(_1108_),
  .S(_1109_)
);

HA_X1 _2187_ (
  .A(result[11]),
  .B(\ext_mult_res[11] ),
  .CO(_1110_),
  .S(_1111_)
);

HA_X1 _2188_ (
  .A(result[12]),
  .B(\ext_mult_res[12] ),
  .CO(_1112_),
  .S(_1113_)
);

HA_X1 _2189_ (
  .A(result[13]),
  .B(\ext_mult_res[13] ),
  .CO(_1114_),
  .S(_1115_)
);

HA_X1 _2190_ (
  .A(result[14]),
  .B(\ext_mult_res[14] ),
  .CO(_1116_),
  .S(_1117_)
);

HA_X1 _2191_ (
  .A(result[15]),
  .B(\ext_mult_res[15] ),
  .CO(_1118_),
  .S(_1119_)
);

HA_X1 _2192_ (
  .A(result[16]),
  .B(\ext_mult_res[16] ),
  .CO(_1120_),
  .S(_1121_)
);

HA_X1 _2193_ (
  .A(result[17]),
  .B(\ext_mult_res[17] ),
  .CO(_1122_),
  .S(_1123_)
);

HA_X1 _2194_ (
  .A(result[18]),
  .B(\ext_mult_res[18] ),
  .CO(_1124_),
  .S(_1125_)
);

HA_X1 _2195_ (
  .A(result[19]),
  .B(\ext_mult_res[18] ),
  .CO(_1126_),
  .S(_1127_)
);

HA_X1 _2196_ (
  .A(result[20]),
  .B(\ext_mult_res[18] ),
  .CO(_1128_),
  .S(_1129_)
);

HA_X1 _2197_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_1132_),
  .S(_1133_)
);

HA_X1 _2198_ (
  .A(_0685_),
  .B(_1132_),
  .CO(_1134_),
  .S(_1135_)
);

HA_X1 _2199_ (
  .A(_0693_),
  .B(_1134_),
  .CO(_1136_),
  .S(_1137_)
);

HA_X1 _2200_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0717_),
  .S(_1140_)
);

HA_X1 _2201_ (
  .A(_1141_),
  .B(_0692_),
  .CO(_1142_),
  .S(_1143_)
);

HA_X1 _2202_ (
  .A(_1143_),
  .B(_1136_),
  .CO(_1144_),
  .S(_1145_)
);

HA_X1 _2203_ (
  .A(_0719_),
  .B(_1142_),
  .CO(_1146_),
  .S(_1147_)
);

HA_X1 _2204_ (
  .A(_1147_),
  .B(_1144_),
  .CO(_1148_),
  .S(_1149_)
);

HA_X1 _2205_ (
  .A(_1150_),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_1152_),
  .S(_1153_)
);

HA_X1 _2206_ (
  .A(_1154_),
  .B(_0718_),
  .CO(_1155_),
  .S(_1156_)
);

HA_X1 _2207_ (
  .A(_1156_),
  .B(_1146_),
  .CO(_1157_),
  .S(_1158_)
);

HA_X1 _2208_ (
  .A(_1158_),
  .B(_1148_),
  .CO(_1159_),
  .S(_1160_)
);

HA_X1 _2209_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_0767_),
  .S(_1162_)
);

HA_X1 _2210_ (
  .A(_1163_),
  .B(_1162_),
  .CO(_0780_),
  .S(_1164_)
);

HA_X1 _2211_ (
  .A(_0782_),
  .B(_1165_),
  .CO(_1166_),
  .S(_1167_)
);

HA_X1 _2212_ (
  .A(_1167_),
  .B(_1168_),
  .CO(_1169_),
  .S(_1170_)
);

HA_X1 _2213_ (
  .A(_1171_),
  .B(_1155_),
  .CO(_1168_),
  .S(_1172_)
);

HA_X1 _2214_ (
  .A(_1170_),
  .B(_1173_),
  .CO(_1174_),
  .S(_1175_)
);

HA_X1 _2215_ (
  .A(_1172_),
  .B(_1157_),
  .CO(_1173_),
  .S(_1176_)
);

HA_X1 _2216_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(_0768_),
  .CO(_0847_),
  .S(_1178_)
);

HA_X1 _2217_ (
  .A(_1179_),
  .B(_0781_),
  .CO(_1180_),
  .S(_1181_)
);

HA_X1 _2218_ (
  .A(_1181_),
  .B(_1166_),
  .CO(_1182_),
  .S(_1183_)
);

HA_X1 _2219_ (
  .A(_1183_),
  .B(_1169_),
  .CO(_1184_),
  .S(_1185_)
);

HA_X1 _2220_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .CO(_1072_),
  .S(_0941_)
);

HA_X1 _2221_ (
  .A(_0814_),
  .B(_0941_),
  .CO(_1186_),
  .S(_1187_)
);

HA_X1 _2222_ (
  .A(_0851_),
  .B(_1180_),
  .CO(_1188_),
  .S(_1189_)
);

HA_X1 _2223_ (
  .A(_1189_),
  .B(_1182_),
  .CO(_1190_),
  .S(_1191_)
);

HA_X1 _2224_ (
  .A(_0875_),
  .B(_1072_),
  .CO(_0910_),
  .S(_1192_)
);

HA_X1 _2225_ (
  .A(_0840_),
  .B(_1192_),
  .CO(_1193_),
  .S(_1194_)
);

HA_X1 _2226_ (
  .A(_0881_),
  .B(_0850_),
  .CO(_1195_),
  .S(_1196_)
);

HA_X1 _2227_ (
  .A(_1196_),
  .B(_1188_),
  .CO(_1197_),
  .S(_1198_)
);

HA_X1 _2228_ (
  .A(_1199_),
  .B(_0918_),
  .CO(_1200_),
  .S(_1201_)
);

HA_X1 _2229_ (
  .A(_1195_),
  .B(_1201_),
  .CO(_1202_),
  .S(_1203_)
);

HA_X1 _2230_ (
  .A(_1204_),
  .B(_1205_),
  .CO(_1206_),
  .S(_1207_)
);

HA_X1 _2231_ (
  .A(_1207_),
  .B(_1200_),
  .CO(_1208_),
  .S(_1209_)
);

HA_X1 _2232_ (
  .A(_1210_),
  .B(_1072_),
  .CO(_1019_),
  .S(_0981_)
);

HA_X1 _2233_ (
  .A(_1211_),
  .B(_0949_),
  .CO(_1212_),
  .S(_1213_)
);

HA_X1 _2234_ (
  .A(_1213_),
  .B(_1206_),
  .CO(_1214_),
  .S(_1215_)
);

HA_X1 _2235_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 ),
  .B(_0874_),
  .CO(_1217_),
  .S(_1218_)
);

HA_X1 _2236_ (
  .A(_0977_),
  .B(_1218_),
  .CO(_1049_),
  .S(_1219_)
);

HA_X1 _2237_ (
  .A(_1021_),
  .B(_1212_),
  .CO(_1220_),
  .S(_1221_)
);

HA_X1 _2238_ (
  .A(_1222_),
  .B(_1216_),
  .CO(_1223_),
  .S(_1224_)
);

HA_X1 _2239_ (
  .A(_0941_),
  .B(_0942_),
  .CO(_1225_),
  .S(_1226_)
);

HA_X1 _2240_ (
  .A(_1226_),
  .B(_1217_),
  .CO(_1077_),
  .S(_1227_)
);

HA_X1 _2241_ (
  .A(_1011_),
  .B(_1227_),
  .CO(_1085_),
  .S(_1228_)
);

HA_X1 _2242_ (
  .A(_1051_),
  .B(_1020_),
  .CO(_1229_),
  .S(_1230_)
);

HA_X1 _2243_ (
  .A(_1074_),
  .B(_1225_),
  .CO(_1231_),
  .S(_1076_)
);

HA_X1 _2244_ (
  .A(_1087_),
  .B(_1050_),
  .CO(_1232_),
  .S(_1233_)
);

HA_X1 _2245_ (
  .A(_1176_),
  .B(_1159_),
  .CO(_1177_),
  .S(_1234_)
);

DFF_X1 \ext_mult_res[0]$_DFFE_PP_  (
  .D(_0000_),
  .CK(clk),
  .Q(\ext_mult_res[0] ),
  .QN(_0675_)
);

DFF_X1 \ext_mult_res[10]$_DFFE_PP_  (
  .D(_0010_),
  .CK(clk),
  .Q(\ext_mult_res[10] ),
  .QN(_0666_)
);

DFF_X1 \ext_mult_res[11]$_DFFE_PP_  (
  .D(_0011_),
  .CK(clk),
  .Q(\ext_mult_res[11] ),
  .QN(_0665_)
);

DFF_X1 \ext_mult_res[12]$_DFFE_PP_  (
  .D(_0012_),
  .CK(clk),
  .Q(\ext_mult_res[12] ),
  .QN(_0664_)
);

DFF_X1 \ext_mult_res[13]$_DFFE_PP_  (
  .D(_0013_),
  .CK(clk),
  .Q(\ext_mult_res[13] ),
  .QN(_0663_)
);

DFF_X1 \ext_mult_res[14]$_DFFE_PP_  (
  .D(_0014_),
  .CK(clk),
  .Q(\ext_mult_res[14] ),
  .QN(_0662_)
);

DFF_X1 \ext_mult_res[15]$_DFFE_PP_  (
  .D(_0015_),
  .CK(clk),
  .Q(\ext_mult_res[15] ),
  .QN(_0661_)
);

DFF_X1 \ext_mult_res[16]$_DFFE_PP_  (
  .D(_0016_),
  .CK(clk),
  .Q(\ext_mult_res[16] ),
  .QN(_0660_)
);

DFF_X1 \ext_mult_res[17]$_DFFE_PP_  (
  .D(_0017_),
  .CK(clk),
  .Q(\ext_mult_res[17] ),
  .QN(_0659_)
);

DFF_X1 \ext_mult_res[1]$_DFFE_PP_  (
  .D(_0001_),
  .CK(clk),
  .Q(\ext_mult_res[1] ),
  .QN(_0677_)
);

DFF_X1 \ext_mult_res[21]$_DFFE_PP_  (
  .D(_0018_),
  .CK(clk),
  .Q(\ext_mult_res[18] ),
  .QN(_0658_)
);

DFF_X1 \ext_mult_res[2]$_DFFE_PP_  (
  .D(_0002_),
  .CK(clk),
  .Q(\ext_mult_res[2] ),
  .QN(_0674_)
);

DFF_X1 \ext_mult_res[3]$_DFFE_PP_  (
  .D(_0003_),
  .CK(clk),
  .Q(\ext_mult_res[3] ),
  .QN(_0673_)
);

DFF_X1 \ext_mult_res[4]$_DFFE_PP_  (
  .D(_0004_),
  .CK(clk),
  .Q(\ext_mult_res[4] ),
  .QN(_0672_)
);

DFF_X1 \ext_mult_res[5]$_DFFE_PP_  (
  .D(_0005_),
  .CK(clk),
  .Q(\ext_mult_res[5] ),
  .QN(_0671_)
);

DFF_X1 \ext_mult_res[6]$_DFFE_PP_  (
  .D(_0006_),
  .CK(clk),
  .Q(\ext_mult_res[6] ),
  .QN(_0670_)
);

DFF_X1 \ext_mult_res[7]$_DFFE_PP_  (
  .D(_0007_),
  .CK(clk),
  .Q(\ext_mult_res[7] ),
  .QN(_0669_)
);

DFF_X1 \ext_mult_res[8]$_DFFE_PP_  (
  .D(_0008_),
  .CK(clk),
  .Q(\ext_mult_res[8] ),
  .QN(_0668_)
);

DFF_X1 \ext_mult_res[9]$_DFFE_PP_  (
  .D(_0009_),
  .CK(clk),
  .Q(\ext_mult_res[9] ),
  .QN(_0667_)
);

DFF_X1 \result[0]$_DFFE_PP_  (
  .D(_0019_),
  .CK(clk),
  .Q(result[0]),
  .QN(_0657_)
);

DFF_X1 \result[10]$_DFFE_PP_  (
  .D(_0029_),
  .CK(clk),
  .Q(result[10]),
  .QN(_0648_)
);

DFF_X1 \result[11]$_DFFE_PP_  (
  .D(_0030_),
  .CK(clk),
  .Q(result[11]),
  .QN(_0647_)
);

DFF_X1 \result[12]$_DFFE_PP_  (
  .D(_0031_),
  .CK(clk),
  .Q(result[12]),
  .QN(_0646_)
);

DFF_X1 \result[13]$_DFFE_PP_  (
  .D(_0032_),
  .CK(clk),
  .Q(result[13]),
  .QN(_0645_)
);

DFF_X1 \result[14]$_DFFE_PP_  (
  .D(_0033_),
  .CK(clk),
  .Q(result[14]),
  .QN(_0644_)
);

DFF_X1 \result[15]$_DFFE_PP_  (
  .D(_0034_),
  .CK(clk),
  .Q(result[15]),
  .QN(_0643_)
);

DFF_X1 \result[16]$_DFFE_PP_  (
  .D(_0035_),
  .CK(clk),
  .Q(result[16]),
  .QN(_0642_)
);

DFF_X1 \result[17]$_DFFE_PP_  (
  .D(_0036_),
  .CK(clk),
  .Q(result[17]),
  .QN(_0641_)
);

DFF_X1 \result[18]$_DFFE_PP_  (
  .D(_0037_),
  .CK(clk),
  .Q(result[18]),
  .QN(_0640_)
);

DFF_X1 \result[19]$_DFFE_PP_  (
  .D(_0038_),
  .CK(clk),
  .Q(result[19]),
  .QN(_0639_)
);

DFF_X1 \result[1]$_DFFE_PP_  (
  .D(_0020_),
  .CK(clk),
  .Q(result[1]),
  .QN(_0676_)
);

DFF_X1 \result[20]$_DFFE_PP_  (
  .D(_0039_),
  .CK(clk),
  .Q(result[20]),
  .QN(_0638_)
);

DFF_X1 \result[21]$_DFFE_PP_  (
  .D(_0040_),
  .CK(clk),
  .Q(result[21]),
  .QN(_0637_)
);

DFF_X1 \result[2]$_DFFE_PP_  (
  .D(_0021_),
  .CK(clk),
  .Q(result[2]),
  .QN(_0656_)
);

DFF_X1 \result[3]$_DFFE_PP_  (
  .D(_0022_),
  .CK(clk),
  .Q(result[3]),
  .QN(_0655_)
);

DFF_X1 \result[4]$_DFFE_PP_  (
  .D(_0023_),
  .CK(clk),
  .Q(result[4]),
  .QN(_0654_)
);

DFF_X1 \result[5]$_DFFE_PP_  (
  .D(_0024_),
  .CK(clk),
  .Q(result[5]),
  .QN(_0653_)
);

DFF_X1 \result[6]$_DFFE_PP_  (
  .D(_0025_),
  .CK(clk),
  .Q(result[6]),
  .QN(_0652_)
);

DFF_X1 \result[7]$_DFFE_PP_  (
  .D(_0026_),
  .CK(clk),
  .Q(result[7]),
  .QN(_0651_)
);

DFF_X1 \result[8]$_DFFE_PP_  (
  .D(_0027_),
  .CK(clk),
  .Q(result[8]),
  .QN(_0650_)
);

DFF_X1 \result[9]$_DFFE_PP_  (
  .D(_0028_),
  .CK(clk),
  .Q(result[9]),
  .QN(_0649_)
);

LOGIC0_X1 \logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974  (
  .Z(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 )
);

LOGIC1_X1 \logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974  (
  .Z(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974 )
);

INV_X1 _1283__reduced (
  .A(_0326_),
  .ZN(_0735_)
);

INV_X1 _1308__reduced (
  .A(_0333_),
  .ZN(_0796_)
);

INV_X1 _1319__reduced (
  .A(_0339_),
  .ZN(_0823_)
);

INV_X1 _1328__reduced (
  .A(_0341_),
  .ZN(_0857_)
);

INV_X1 _1337__reduced (
  .A(_0354_),
  .ZN(_0886_)
);

INV_X1 _1345__reduced (
  .A(_0355_),
  .ZN(_0921_)
);

INV_X1 _1353__reduced (
  .A(_0348_),
  .ZN(_0959_)
);

INV_X1 _1359__reduced (
  .A(din[7]),
  .ZN(_0993_)
);

NOR2_X1 _1473__reduced (
  .A1(_0370_),
  .A2(_0372_),
  .ZN(_0000_)
);

INV_X1 _1634__reduced (
  .A(_0993_),
  .ZN(_0516_)
);

INV_X1 _1636__reduced (
  .A(_0516_),
  .ZN(_0518_)
);

NAND2_X1 _1638__reduced (
  .A1(_0516_),
  .A2(_0358_),
  .ZN(_0520_)
);

NAND2_X1 _1643__reduced (
  .A1(_0516_),
  .A2(_0524_),
  .ZN(_0525_)
);

NAND2_X1 _1662__reduced (
  .A1(_0540_),
  .A2(_0541_),
  .ZN(_0544_)
);

INV_X1 _1663__reduced (
  .A(_0544_),
  .ZN(_0545_)
);

NAND2_X1 _1667__reduced (
  .A1(_0544_),
  .A2(_0546_),
  .ZN(_0549_)
);
endmodule //$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974

module jpeg_rzs_clone_498(input clk, input ena, input rst, input deni, input dci,
 input [3:0] rleni, input [3:0] sizei, input [11:0] ampi, output deno, output dco, output [3:0] rleno,
 output [3:0] sizeo, output [11:0] ampo);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire \amp[0] ;
wire \amp[10] ;
wire \amp[11] ;
wire \amp[1] ;
wire \amp[2] ;
wire \amp[3] ;
wire \amp[4] ;
wire \amp[5] ;
wire \amp[6] ;
wire \amp[7] ;
wire \amp[8] ;
wire \amp[9] ;
wire dc;
wire den;
wire \rlen[0] ;
wire \rlen[1] ;
wire \rlen[2] ;
wire \rlen[3] ;
wire \size[0] ;
wire \size[1] ;
wire \size[2] ;
wire \size[3] ;
wire state;

NAND2_X1 _120_ (
  .A1(rleni[1]),
  .A2(rleni[0]),
  .ZN(_045_)
);

NAND2_X1 _121_ (
  .A1(rleni[3]),
  .A2(rleni[2]),
  .ZN(_046_)
);

NOR2_X1 _122_ (
  .A1(_045_),
  .A2(_046_),
  .ZN(_047_)
);

NOR2_X1 _123_ (
  .A1(sizei[1]),
  .A2(sizei[0]),
  .ZN(_048_)
);

NOR2_X1 _124_ (
  .A1(sizei[3]),
  .A2(sizei[2]),
  .ZN(_049_)
);

NAND3_X1 _125_ (
  .A1(_047_),
  .A2(_048_),
  .A3(_049_),
  .ZN(_050_)
);

BUF_X4 _126_ (
  .A(ena),
  .Z(_051_)
);

NAND2_X4 _127_ (
  .A1(deni),
  .A2(_051_),
  .ZN(_052_)
);

BUF_X8 _128_ (
  .A(_052_),
  .Z(_053_)
);

INV_X1 _129_ (
  .A(_053_),
  .ZN(_054_)
);

NAND2_X1 _130_ (
  .A1(_050_),
  .A2(_054_),
  .ZN(_055_)
);

INV_X1 _131_ (
  .A(state),
  .ZN(_056_)
);

NAND2_X1 _132_ (
  .A1(_056_),
  .A2(_051_),
  .ZN(_057_)
);

NAND3_X1 _133_ (
  .A1(_057_),
  .A2(_053_),
  .A3(den),
  .ZN(_058_)
);

NAND2_X1 _134_ (
  .A1(_055_),
  .A2(_058_),
  .ZN(_000_)
);

NOR2_X1 _135_ (
  .A1(_052_),
  .A2(_056_),
  .ZN(_059_)
);

NOR2_X1 _136_ (
  .A1(rleni[1]),
  .A2(rleni[0]),
  .ZN(_060_)
);

NOR2_X1 _137_ (
  .A1(rleni[3]),
  .A2(rleni[2]),
  .ZN(_061_)
);

INV_X1 _138_ (
  .A(dci),
  .ZN(_062_)
);

NAND3_X1 _139_ (
  .A1(_060_),
  .A2(_061_),
  .A3(_062_),
  .ZN(_063_)
);

NAND2_X1 _140_ (
  .A1(_048_),
  .A2(_049_),
  .ZN(_064_)
);

OAI21_X1 _141_ (
  .A(_059_),
  .B1(_063_),
  .B2(_064_),
  .ZN(_065_)
);

INV_X1 _142_ (
  .A(den),
  .ZN(_066_)
);

INV_X1 _143_ (
  .A(deno),
  .ZN(_067_)
);

OAI22_X1 _144_ (
  .A1(_057_),
  .A2(_066_),
  .B1(_067_),
  .B2(_051_),
  .ZN(_068_)
);

INV_X1 _145_ (
  .A(_068_),
  .ZN(_069_)
);

NAND2_X1 _146_ (
  .A1(_065_),
  .A2(_069_),
  .ZN(_001_)
);

BUF_X4 _147_ (
  .A(_051_),
  .Z(_070_)
);

NOR2_X1 _148_ (
  .A1(_070_),
  .A2(dc),
  .ZN(_071_)
);

AOI21_X1 _149_ (
  .A(_071_),
  .B1(_062_),
  .B2(_070_),
  .ZN(_002_)
);

BUF_X4 _150_ (
  .A(_051_),
  .Z(_072_)
);

MUX2_X1 _151_ (
  .A(rleno[0]),
  .B(\rlen[0] ),
  .S(_072_),
  .Z(_003_)
);

MUX2_X1 _152_ (
  .A(rleno[1]),
  .B(\rlen[1] ),
  .S(_070_),
  .Z(_004_)
);

MUX2_X1 _153_ (
  .A(rleno[2]),
  .B(\rlen[2] ),
  .S(_072_),
  .Z(_005_)
);

MUX2_X1 _154_ (
  .A(rleno[3]),
  .B(\rlen[3] ),
  .S(_070_),
  .Z(_006_)
);

MUX2_X1 _155_ (
  .A(sizeo[0]),
  .B(\size[0] ),
  .S(_072_),
  .Z(_007_)
);

MUX2_X1 _156_ (
  .A(sizeo[1]),
  .B(\size[1] ),
  .S(_051_),
  .Z(_008_)
);

MUX2_X1 _157_ (
  .A(sizeo[2]),
  .B(\size[2] ),
  .S(_051_),
  .Z(_009_)
);

MUX2_X1 _158_ (
  .A(sizeo[3]),
  .B(\size[3] ),
  .S(_070_),
  .Z(_010_)
);

MUX2_X1 _159_ (
  .A(ampo[0]),
  .B(\amp[0] ),
  .S(_072_),
  .Z(_011_)
);

MUX2_X1 _160_ (
  .A(ampo[1]),
  .B(\amp[1] ),
  .S(_072_),
  .Z(_012_)
);

MUX2_X1 _161_ (
  .A(ampo[2]),
  .B(\amp[2] ),
  .S(_070_),
  .Z(_013_)
);

MUX2_X1 _162_ (
  .A(ampo[3]),
  .B(\amp[3] ),
  .S(_072_),
  .Z(_014_)
);

MUX2_X1 _163_ (
  .A(ampo[4]),
  .B(\amp[4] ),
  .S(_070_),
  .Z(_015_)
);

MUX2_X1 _164_ (
  .A(ampo[5]),
  .B(\amp[5] ),
  .S(_072_),
  .Z(_016_)
);

MUX2_X1 _165_ (
  .A(ampo[6]),
  .B(\amp[6] ),
  .S(_070_),
  .Z(_017_)
);

MUX2_X1 _166_ (
  .A(ampo[7]),
  .B(\amp[7] ),
  .S(_072_),
  .Z(_018_)
);

MUX2_X1 _167_ (
  .A(ampo[8]),
  .B(\amp[8] ),
  .S(_072_),
  .Z(_019_)
);

MUX2_X1 _168_ (
  .A(ampo[9]),
  .B(\amp[9] ),
  .S(_070_),
  .Z(_020_)
);

MUX2_X1 _169_ (
  .A(ampo[10]),
  .B(\amp[10] ),
  .S(_072_),
  .Z(_021_)
);

MUX2_X1 _170_ (
  .A(ampo[11]),
  .B(\amp[11] ),
  .S(_070_),
  .Z(_022_)
);

MUX2_X1 _171_ (
  .A(dco),
  .B(dc),
  .S(_051_),
  .Z(_023_)
);

MUX2_X1 _172_ (
  .A(sizei[0]),
  .B(\size[0] ),
  .S(_053_),
  .Z(_024_)
);

BUF_X8 _173_ (
  .A(_052_),
  .Z(_073_)
);

MUX2_X1 _174_ (
  .A(sizei[1]),
  .B(\size[1] ),
  .S(_073_),
  .Z(_025_)
);

MUX2_X1 _175_ (
  .A(sizei[2]),
  .B(\size[2] ),
  .S(_053_),
  .Z(_026_)
);

MUX2_X1 _176_ (
  .A(sizei[3]),
  .B(\size[3] ),
  .S(_053_),
  .Z(_027_)
);

MUX2_X1 _177_ (
  .A(rleni[0]),
  .B(\rlen[0] ),
  .S(_053_),
  .Z(_028_)
);

MUX2_X1 _178_ (
  .A(rleni[1]),
  .B(\rlen[1] ),
  .S(_053_),
  .Z(_029_)
);

MUX2_X1 _179_ (
  .A(rleni[2]),
  .B(\rlen[2] ),
  .S(_053_),
  .Z(_030_)
);

MUX2_X1 _180_ (
  .A(rleni[3]),
  .B(\rlen[3] ),
  .S(_073_),
  .Z(_031_)
);

MUX2_X1 _181_ (
  .A(ampi[0]),
  .B(\amp[0] ),
  .S(_073_),
  .Z(_032_)
);

MUX2_X1 _182_ (
  .A(ampi[1]),
  .B(\amp[1] ),
  .S(_073_),
  .Z(_033_)
);

MUX2_X1 _183_ (
  .A(ampi[2]),
  .B(\amp[2] ),
  .S(_073_),
  .Z(_034_)
);

MUX2_X1 _184_ (
  .A(ampi[3]),
  .B(\amp[3] ),
  .S(_052_),
  .Z(_035_)
);

MUX2_X1 _185_ (
  .A(ampi[4]),
  .B(\amp[4] ),
  .S(_073_),
  .Z(_036_)
);

MUX2_X1 _186_ (
  .A(ampi[5]),
  .B(\amp[5] ),
  .S(_073_),
  .Z(_037_)
);

MUX2_X1 _187_ (
  .A(ampi[6]),
  .B(\amp[6] ),
  .S(_073_),
  .Z(_038_)
);

MUX2_X1 _188_ (
  .A(ampi[7]),
  .B(\amp[7] ),
  .S(_073_),
  .Z(_039_)
);

MUX2_X1 _189_ (
  .A(ampi[8]),
  .B(\amp[8] ),
  .S(_073_),
  .Z(_040_)
);

MUX2_X1 _190_ (
  .A(ampi[9]),
  .B(\amp[9] ),
  .S(_052_),
  .Z(_041_)
);

MUX2_X1 _191_ (
  .A(ampi[10]),
  .B(\amp[10] ),
  .S(_052_),
  .Z(_042_)
);

NAND2_X1 _193_ (
  .A1(_053_),
  .A2(state),
  .ZN(_074_)
);

OAI21_X1 _194_ (
  .A(_074_),
  .B1(_050_),
  .B2(_053_),
  .ZN(_044_)
);

DFF_X1 \amp[0]$_DFFE_PP_  (
  .D(_032_),
  .CK(clk),
  .Q(\amp[0] ),
  .QN(_087_)
);

DFF_X1 \amp[10]$_DFFE_PP_  (
  .D(_042_),
  .CK(clk),
  .Q(\amp[10] ),
  .QN(_077_)
);

DFF_X1 \amp[11]$_DFFE_PP_  (
  .D(_043_),
  .CK(clk),
  .Q(\amp[11] ),
  .QN(_076_)
);

DFF_X1 \amp[1]$_DFFE_PP_  (
  .D(_033_),
  .CK(clk),
  .Q(\amp[1] ),
  .QN(_086_)
);

DFF_X1 \amp[2]$_DFFE_PP_  (
  .D(_034_),
  .CK(clk),
  .Q(\amp[2] ),
  .QN(_085_)
);

DFF_X1 \amp[3]$_DFFE_PP_  (
  .D(_035_),
  .CK(clk),
  .Q(\amp[3] ),
  .QN(_084_)
);

DFF_X1 \amp[4]$_DFFE_PP_  (
  .D(_036_),
  .CK(clk),
  .Q(\amp[4] ),
  .QN(_083_)
);

DFF_X1 \amp[5]$_DFFE_PP_  (
  .D(_037_),
  .CK(clk),
  .Q(\amp[5] ),
  .QN(_082_)
);

DFF_X1 \amp[6]$_DFFE_PP_  (
  .D(_038_),
  .CK(clk),
  .Q(\amp[6] ),
  .QN(_081_)
);

DFF_X1 \amp[7]$_DFFE_PP_  (
  .D(_039_),
  .CK(clk),
  .Q(\amp[7] ),
  .QN(_080_)
);

DFF_X1 \amp[8]$_DFFE_PP_  (
  .D(_040_),
  .CK(clk),
  .Q(\amp[8] ),
  .QN(_079_)
);

DFF_X1 \amp[9]$_DFFE_PP_  (
  .D(_041_),
  .CK(clk),
  .Q(\amp[9] ),
  .QN(_078_)
);

DFF_X1 \ampo[0]$_DFFE_PP_  (
  .D(_011_),
  .CK(clk),
  .Q(ampo[0]),
  .QN(_108_)
);

DFF_X1 \ampo[10]$_DFFE_PP_  (
  .D(_021_),
  .CK(clk),
  .Q(ampo[10]),
  .QN(_098_)
);

DFF_X1 \ampo[11]$_DFFE_PP_  (
  .D(_022_),
  .CK(clk),
  .Q(ampo[11]),
  .QN(_097_)
);

DFF_X1 \ampo[1]$_DFFE_PP_  (
  .D(_012_),
  .CK(clk),
  .Q(ampo[1]),
  .QN(_107_)
);

DFF_X1 \ampo[2]$_DFFE_PP_  (
  .D(_013_),
  .CK(clk),
  .Q(ampo[2]),
  .QN(_106_)
);

DFF_X1 \ampo[3]$_DFFE_PP_  (
  .D(_014_),
  .CK(clk),
  .Q(ampo[3]),
  .QN(_105_)
);

DFF_X1 \ampo[4]$_DFFE_PP_  (
  .D(_015_),
  .CK(clk),
  .Q(ampo[4]),
  .QN(_104_)
);

DFF_X1 \ampo[5]$_DFFE_PP_  (
  .D(_016_),
  .CK(clk),
  .Q(ampo[5]),
  .QN(_103_)
);

DFF_X1 \ampo[6]$_DFFE_PP_  (
  .D(_017_),
  .CK(clk),
  .Q(ampo[6]),
  .QN(_102_)
);

DFF_X1 \ampo[7]$_DFFE_PP_  (
  .D(_018_),
  .CK(clk),
  .Q(ampo[7]),
  .QN(_101_)
);

DFF_X1 \ampo[8]$_DFFE_PP_  (
  .D(_019_),
  .CK(clk),
  .Q(ampo[8]),
  .QN(_100_)
);

DFF_X1 \ampo[9]$_DFFE_PP_  (
  .D(_020_),
  .CK(clk),
  .Q(ampo[9]),
  .QN(_099_)
);

DFF_X1 dc$_DFFE_PP_ (
  .D(_002_),
  .CK(clk),
  .Q(dc),
  .QN(_117_)
);

DFF_X1 dco$_DFFE_PP_ (
  .D(_023_),
  .CK(clk),
  .Q(dco),
  .QN(_096_)
);

DFFR_X1 den$_DFFE_PN0P_ (
  .D(_000_),
  .RN(rst),
  .CK(clk),
  .Q(den),
  .QN(_119_)
);

DFFR_X1 deno$_DFFE_PN0P_ (
  .D(_001_),
  .RN(rst),
  .CK(clk),
  .Q(deno),
  .QN(_118_)
);

DFF_X1 \rlen[0]$_DFFE_PP_  (
  .D(_028_),
  .CK(clk),
  .Q(\rlen[0] ),
  .QN(_091_)
);

DFF_X1 \rlen[1]$_DFFE_PP_  (
  .D(_029_),
  .CK(clk),
  .Q(\rlen[1] ),
  .QN(_090_)
);

DFF_X1 \rlen[2]$_DFFE_PP_  (
  .D(_030_),
  .CK(clk),
  .Q(\rlen[2] ),
  .QN(_089_)
);

DFF_X1 \rlen[3]$_DFFE_PP_  (
  .D(_031_),
  .CK(clk),
  .Q(\rlen[3] ),
  .QN(_088_)
);

DFF_X1 \rleno[0]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(rleno[0]),
  .QN(_116_)
);

DFF_X1 \rleno[1]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(rleno[1]),
  .QN(_115_)
);

DFF_X1 \rleno[2]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(rleno[2]),
  .QN(_114_)
);

DFF_X1 \rleno[3]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(rleno[3]),
  .QN(_113_)
);

DFF_X1 \size[0]$_DFFE_PP_  (
  .D(_024_),
  .CK(clk),
  .Q(\size[0] ),
  .QN(_095_)
);

DFF_X1 \size[1]$_DFFE_PP_  (
  .D(_025_),
  .CK(clk),
  .Q(\size[1] ),
  .QN(_094_)
);

DFF_X1 \size[2]$_DFFE_PP_  (
  .D(_026_),
  .CK(clk),
  .Q(\size[2] ),
  .QN(_093_)
);

DFF_X1 \size[3]$_DFFE_PP_  (
  .D(_027_),
  .CK(clk),
  .Q(\size[3] ),
  .QN(_092_)
);

DFF_X1 \sizeo[0]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(sizeo[0]),
  .QN(_112_)
);

DFF_X1 \sizeo[1]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(sizeo[1]),
  .QN(_111_)
);

DFF_X1 \sizeo[2]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(sizeo[2]),
  .QN(_110_)
);

DFF_X1 \sizeo[3]$_DFFE_PP_  (
  .D(_010_),
  .CK(clk),
  .Q(sizeo[3]),
  .QN(_109_)
);

DFFR_X1 state$_DFFE_PN0P_ (
  .D(_044_),
  .RN(rst),
  .CK(clk),
  .Q(state),
  .QN(_075_)
);

AND2_X1 _192__reduced (
  .A1(\amp[11] ),
  .A2(_052_),
  .ZN(_043_)
);
endmodule //jpeg_rzs_clone_498

module zigzag(input clk, input ena, input dstrb, input [11:0] din_00, input [11:0] din_01,
 input [11:0] din_02, input [11:0] din_03, input [11:0] din_04, input [11:0] din_05, input [11:0] din_06,
 input [11:0] din_07, input [11:0] din_10, input [11:0] din_11, input [11:0] din_12, input [11:0] din_13,
 input [11:0] din_14, input [11:0] din_15, input [11:0] din_16, input [11:0] din_17, input [11:0] din_20,
 input [11:0] din_21, input [11:0] din_22, input [11:0] din_23, input [11:0] din_24, input [11:0] din_25,
 input [11:0] din_26, input [11:0] din_27, input [11:0] din_30, input [11:0] din_31, input [11:0] din_32,
 input [11:0] din_33, input [11:0] din_34, input [11:0] din_35, input [11:0] din_36, input [11:0] din_37,
 input [11:0] din_40, input [11:0] din_41, input [11:0] din_42, input [11:0] din_43, input [11:0] din_44,
 input [11:0] din_45, input [11:0] din_46, input [11:0] din_47, input [11:0] din_50, input [11:0] din_51,
 input [11:0] din_52, input [11:0] din_53, input [11:0] din_54, input [11:0] din_55, input [11:0] din_56,
 input [11:0] din_57, input [11:0] din_60, input [11:0] din_61, input [11:0] din_62, input [11:0] din_63,
 input [11:0] din_64, input [11:0] din_65, input [11:0] din_66, input [11:0] din_67, input [11:0] din_70,
 input [11:0] din_71, input [11:0] din_72, input [11:0] din_73, input [11:0] din_74, input [11:0] din_75,
 input [11:0] din_76, input [11:0] din_77, output [11:0] dout, output douten);
wire _00000_;
wire _00001_;
wire _00002_;
wire _00003_;
wire _00004_;
wire _00005_;
wire _00006_;
wire _00007_;
wire _00008_;
wire _00009_;
wire _00010_;
wire _00011_;
wire _00012_;
wire _00013_;
wire _00014_;
wire _00015_;
wire _00016_;
wire _00017_;
wire _00018_;
wire _00019_;
wire _00020_;
wire _00021_;
wire _00022_;
wire _00023_;
wire _00024_;
wire _00025_;
wire _00026_;
wire _00027_;
wire _00028_;
wire _00029_;
wire _00030_;
wire _00031_;
wire _00032_;
wire _00033_;
wire _00034_;
wire _00035_;
wire _00036_;
wire _00037_;
wire _00038_;
wire _00039_;
wire _00040_;
wire _00041_;
wire _00042_;
wire _00043_;
wire _00044_;
wire _00045_;
wire _00046_;
wire _00047_;
wire _00048_;
wire _00049_;
wire _00050_;
wire _00051_;
wire _00052_;
wire _00053_;
wire _00054_;
wire _00055_;
wire _00056_;
wire _00057_;
wire _00058_;
wire _00059_;
wire _00060_;
wire _00061_;
wire _00062_;
wire _00063_;
wire _00064_;
wire _00065_;
wire _00066_;
wire _00067_;
wire _00068_;
wire _00069_;
wire _00070_;
wire _00071_;
wire _00072_;
wire _00073_;
wire _00074_;
wire _00075_;
wire _00076_;
wire _00077_;
wire _00078_;
wire _00079_;
wire _00080_;
wire _00081_;
wire _00082_;
wire _00083_;
wire _00084_;
wire _00085_;
wire _00086_;
wire _00087_;
wire _00088_;
wire _00089_;
wire _00090_;
wire _00091_;
wire _00092_;
wire _00093_;
wire _00094_;
wire _00095_;
wire _00096_;
wire _00097_;
wire _00098_;
wire _00099_;
wire _00100_;
wire _00101_;
wire _00102_;
wire _00103_;
wire _00104_;
wire _00105_;
wire _00106_;
wire _00107_;
wire _00108_;
wire _00109_;
wire _00110_;
wire _00111_;
wire _00112_;
wire _00113_;
wire _00114_;
wire _00115_;
wire _00116_;
wire _00117_;
wire _00118_;
wire _00119_;
wire _00120_;
wire _00121_;
wire _00122_;
wire _00123_;
wire _00124_;
wire _00125_;
wire _00126_;
wire _00127_;
wire _00128_;
wire _00129_;
wire _00130_;
wire _00131_;
wire _00132_;
wire _00133_;
wire _00134_;
wire _00135_;
wire _00136_;
wire _00137_;
wire _00138_;
wire _00139_;
wire _00140_;
wire _00141_;
wire _00142_;
wire _00143_;
wire _00144_;
wire _00145_;
wire _00146_;
wire _00147_;
wire _00148_;
wire _00149_;
wire _00150_;
wire _00151_;
wire _00152_;
wire _00153_;
wire _00154_;
wire _00155_;
wire _00156_;
wire _00157_;
wire _00158_;
wire _00159_;
wire _00160_;
wire _00161_;
wire _00162_;
wire _00163_;
wire _00164_;
wire _00165_;
wire _00166_;
wire _00167_;
wire _00168_;
wire _00169_;
wire _00170_;
wire _00171_;
wire _00172_;
wire _00173_;
wire _00174_;
wire _00175_;
wire _00176_;
wire _00177_;
wire _00178_;
wire _00179_;
wire _00180_;
wire _00181_;
wire _00182_;
wire _00183_;
wire _00184_;
wire _00185_;
wire _00186_;
wire _00187_;
wire _00188_;
wire _00189_;
wire _00190_;
wire _00191_;
wire _00192_;
wire _00193_;
wire _00194_;
wire _00195_;
wire _00196_;
wire _00197_;
wire _00198_;
wire _00199_;
wire _00200_;
wire _00201_;
wire _00202_;
wire _00203_;
wire _00204_;
wire _00205_;
wire _00206_;
wire _00207_;
wire _00208_;
wire _00209_;
wire _00210_;
wire _00211_;
wire _00212_;
wire _00213_;
wire _00214_;
wire _00215_;
wire _00216_;
wire _00217_;
wire _00218_;
wire _00219_;
wire _00220_;
wire _00221_;
wire _00222_;
wire _00223_;
wire _00224_;
wire _00225_;
wire _00226_;
wire _00227_;
wire _00228_;
wire _00229_;
wire _00230_;
wire _00231_;
wire _00232_;
wire _00233_;
wire _00234_;
wire _00235_;
wire _00236_;
wire _00237_;
wire _00238_;
wire _00239_;
wire _00240_;
wire _00241_;
wire _00242_;
wire _00243_;
wire _00244_;
wire _00245_;
wire _00246_;
wire _00247_;
wire _00248_;
wire _00249_;
wire _00250_;
wire _00251_;
wire _00252_;
wire _00253_;
wire _00254_;
wire _00255_;
wire _00256_;
wire _00257_;
wire _00258_;
wire _00259_;
wire _00260_;
wire _00261_;
wire _00262_;
wire _00263_;
wire _00264_;
wire _00265_;
wire _00266_;
wire _00267_;
wire _00268_;
wire _00269_;
wire _00270_;
wire _00271_;
wire _00272_;
wire _00273_;
wire _00274_;
wire _00275_;
wire _00276_;
wire _00277_;
wire _00278_;
wire _00279_;
wire _00280_;
wire _00281_;
wire _00282_;
wire _00283_;
wire _00284_;
wire _00285_;
wire _00286_;
wire _00287_;
wire _00288_;
wire _00289_;
wire _00290_;
wire _00291_;
wire _00292_;
wire _00293_;
wire _00294_;
wire _00295_;
wire _00296_;
wire _00297_;
wire _00298_;
wire _00299_;
wire _00300_;
wire _00301_;
wire _00302_;
wire _00303_;
wire _00304_;
wire _00305_;
wire _00306_;
wire _00307_;
wire _00308_;
wire _00309_;
wire _00310_;
wire _00311_;
wire _00312_;
wire _00313_;
wire _00314_;
wire _00315_;
wire _00316_;
wire _00317_;
wire _00318_;
wire _00319_;
wire _00320_;
wire _00321_;
wire _00322_;
wire _00323_;
wire _00324_;
wire _00325_;
wire _00326_;
wire _00327_;
wire _00328_;
wire _00329_;
wire _00330_;
wire _00331_;
wire _00332_;
wire _00333_;
wire _00334_;
wire _00335_;
wire _00336_;
wire _00337_;
wire _00338_;
wire _00339_;
wire _00340_;
wire _00341_;
wire _00342_;
wire _00343_;
wire _00344_;
wire _00345_;
wire _00346_;
wire _00347_;
wire _00348_;
wire _00349_;
wire _00350_;
wire _00351_;
wire _00352_;
wire _00353_;
wire _00354_;
wire _00355_;
wire _00356_;
wire _00357_;
wire _00358_;
wire _00359_;
wire _00360_;
wire _00361_;
wire _00362_;
wire _00363_;
wire _00364_;
wire _00365_;
wire _00366_;
wire _00367_;
wire _00368_;
wire _00369_;
wire _00370_;
wire _00371_;
wire _00372_;
wire _00373_;
wire _00374_;
wire _00375_;
wire _00376_;
wire _00377_;
wire _00378_;
wire _00379_;
wire _00380_;
wire _00381_;
wire _00382_;
wire _00383_;
wire _00384_;
wire _00385_;
wire _00386_;
wire _00387_;
wire _00388_;
wire _00389_;
wire _00390_;
wire _00391_;
wire _00392_;
wire _00393_;
wire _00394_;
wire _00395_;
wire _00396_;
wire _00397_;
wire _00398_;
wire _00399_;
wire _00400_;
wire _00401_;
wire _00402_;
wire _00403_;
wire _00404_;
wire _00405_;
wire _00406_;
wire _00407_;
wire _00408_;
wire _00409_;
wire _00410_;
wire _00411_;
wire _00412_;
wire _00413_;
wire _00414_;
wire _00415_;
wire _00416_;
wire _00417_;
wire _00418_;
wire _00419_;
wire _00420_;
wire _00421_;
wire _00422_;
wire _00423_;
wire _00424_;
wire _00425_;
wire _00426_;
wire _00427_;
wire _00428_;
wire _00429_;
wire _00430_;
wire _00431_;
wire _00432_;
wire _00433_;
wire _00434_;
wire _00435_;
wire _00436_;
wire _00437_;
wire _00438_;
wire _00439_;
wire _00440_;
wire _00441_;
wire _00442_;
wire _00443_;
wire _00444_;
wire _00445_;
wire _00446_;
wire _00447_;
wire _00448_;
wire _00449_;
wire _00450_;
wire _00451_;
wire _00452_;
wire _00453_;
wire _00454_;
wire _00455_;
wire _00456_;
wire _00457_;
wire _00458_;
wire _00459_;
wire _00460_;
wire _00461_;
wire _00462_;
wire _00463_;
wire _00464_;
wire _00465_;
wire _00466_;
wire _00467_;
wire _00468_;
wire _00469_;
wire _00470_;
wire _00471_;
wire _00472_;
wire _00473_;
wire _00474_;
wire _00475_;
wire _00476_;
wire _00477_;
wire _00478_;
wire _00479_;
wire _00480_;
wire _00481_;
wire _00482_;
wire _00483_;
wire _00484_;
wire _00485_;
wire _00486_;
wire _00487_;
wire _00488_;
wire _00489_;
wire _00490_;
wire _00491_;
wire _00492_;
wire _00493_;
wire _00494_;
wire _00495_;
wire _00496_;
wire _00497_;
wire _00498_;
wire _00499_;
wire _00500_;
wire _00501_;
wire _00502_;
wire _00503_;
wire _00504_;
wire _00505_;
wire _00506_;
wire _00507_;
wire _00508_;
wire _00509_;
wire _00510_;
wire _00511_;
wire _00512_;
wire _00513_;
wire _00514_;
wire _00515_;
wire _00516_;
wire _00517_;
wire _00518_;
wire _00519_;
wire _00520_;
wire _00521_;
wire _00522_;
wire _00523_;
wire _00524_;
wire _00525_;
wire _00526_;
wire _00527_;
wire _00528_;
wire _00529_;
wire _00530_;
wire _00531_;
wire _00532_;
wire _00533_;
wire _00534_;
wire _00535_;
wire _00536_;
wire _00537_;
wire _00538_;
wire _00539_;
wire _00540_;
wire _00541_;
wire _00542_;
wire _00543_;
wire _00544_;
wire _00545_;
wire _00546_;
wire _00547_;
wire _00548_;
wire _00549_;
wire _00550_;
wire _00551_;
wire _00552_;
wire _00553_;
wire _00554_;
wire _00555_;
wire _00556_;
wire _00557_;
wire _00558_;
wire _00559_;
wire _00560_;
wire _00561_;
wire _00562_;
wire _00563_;
wire _00564_;
wire _00565_;
wire _00566_;
wire _00567_;
wire _00568_;
wire _00569_;
wire _00570_;
wire _00571_;
wire _00572_;
wire _00573_;
wire _00574_;
wire _00575_;
wire _00576_;
wire _00577_;
wire _00578_;
wire _00579_;
wire _00580_;
wire _00581_;
wire _00582_;
wire _00583_;
wire _00584_;
wire _00585_;
wire _00586_;
wire _00587_;
wire _00588_;
wire _00589_;
wire _00590_;
wire _00591_;
wire _00592_;
wire _00593_;
wire _00594_;
wire _00595_;
wire _00596_;
wire _00597_;
wire _00598_;
wire _00599_;
wire _00600_;
wire _00601_;
wire _00602_;
wire _00603_;
wire _00604_;
wire _00605_;
wire _00606_;
wire _00607_;
wire _00608_;
wire _00609_;
wire _00610_;
wire _00611_;
wire _00612_;
wire _00613_;
wire _00614_;
wire _00615_;
wire _00616_;
wire _00617_;
wire _00618_;
wire _00619_;
wire _00620_;
wire _00621_;
wire _00622_;
wire _00623_;
wire _00624_;
wire _00625_;
wire _00626_;
wire _00627_;
wire _00628_;
wire _00629_;
wire _00630_;
wire _00631_;
wire _00632_;
wire _00633_;
wire _00634_;
wire _00635_;
wire _00636_;
wire _00637_;
wire _00638_;
wire _00639_;
wire _00640_;
wire _00641_;
wire _00642_;
wire _00643_;
wire _00644_;
wire _00645_;
wire _00646_;
wire _00647_;
wire _00648_;
wire _00649_;
wire _00650_;
wire _00651_;
wire _00652_;
wire _00653_;
wire _00654_;
wire _00655_;
wire _00656_;
wire _00657_;
wire _00658_;
wire _00659_;
wire _00660_;
wire _00661_;
wire _00662_;
wire _00663_;
wire _00664_;
wire _00665_;
wire _00666_;
wire _00667_;
wire _00668_;
wire _00669_;
wire _00670_;
wire _00671_;
wire _00672_;
wire _00673_;
wire _00674_;
wire _00675_;
wire _00676_;
wire _00677_;
wire _00678_;
wire _00679_;
wire _00680_;
wire _00681_;
wire _00682_;
wire _00683_;
wire _00684_;
wire _00685_;
wire _00686_;
wire _00687_;
wire _00688_;
wire _00689_;
wire _00690_;
wire _00691_;
wire _00692_;
wire _00693_;
wire _00694_;
wire _00695_;
wire _00696_;
wire _00697_;
wire _00698_;
wire _00699_;
wire _00700_;
wire _00701_;
wire _00702_;
wire _00703_;
wire _00704_;
wire _00705_;
wire _00706_;
wire _00707_;
wire _00708_;
wire _00709_;
wire _00710_;
wire _00711_;
wire _00712_;
wire _00713_;
wire _00714_;
wire _00715_;
wire _00716_;
wire _00717_;
wire _00718_;
wire _00719_;
wire _00720_;
wire _00721_;
wire _00722_;
wire _00723_;
wire _00724_;
wire _00725_;
wire _00726_;
wire _00727_;
wire _00728_;
wire _00729_;
wire _00730_;
wire _00731_;
wire _00732_;
wire _00733_;
wire _00734_;
wire _00735_;
wire _00736_;
wire _00737_;
wire _00738_;
wire _00739_;
wire _00740_;
wire _00741_;
wire _00742_;
wire _00743_;
wire _00744_;
wire _00745_;
wire _00746_;
wire _00747_;
wire _00748_;
wire _00749_;
wire _00750_;
wire _00751_;
wire _00752_;
wire _00753_;
wire _00754_;
wire _00755_;
wire _00756_;
wire _00757_;
wire _00758_;
wire _00759_;
wire _00760_;
wire _00761_;
wire _00762_;
wire _00763_;
wire _00764_;
wire _00765_;
wire _00766_;
wire _00767_;
wire _00768_;
wire _00769_;
wire _00770_;
wire _00771_;
wire _00772_;
wire _00773_;
wire _00774_;
wire _00775_;
wire _00776_;
wire _00777_;
wire _00778_;
wire _00779_;
wire _00780_;
wire _00781_;
wire _00782_;
wire _00783_;
wire _00784_;
wire _00785_;
wire _00786_;
wire _00787_;
wire _00788_;
wire _00789_;
wire _00790_;
wire _00791_;
wire _00792_;
wire _00793_;
wire _00794_;
wire _00795_;
wire _00796_;
wire _00797_;
wire _00798_;
wire _00799_;
wire _00800_;
wire _00801_;
wire _00802_;
wire _00803_;
wire _00804_;
wire _00805_;
wire _00806_;
wire _00807_;
wire _00808_;
wire _00809_;
wire _00810_;
wire _00811_;
wire _00812_;
wire _00813_;
wire _00814_;
wire _00815_;
wire _00816_;
wire _00817_;
wire _00818_;
wire _00819_;
wire _00820_;
wire _00821_;
wire _00822_;
wire _00823_;
wire _00824_;
wire _00825_;
wire _00826_;
wire _00827_;
wire _00828_;
wire _00829_;
wire _00830_;
wire _00831_;
wire _00832_;
wire _00833_;
wire _00834_;
wire _00835_;
wire _00836_;
wire _00837_;
wire _00838_;
wire _00839_;
wire _00840_;
wire _00841_;
wire _00842_;
wire _00843_;
wire _00844_;
wire _00845_;
wire _00846_;
wire _00847_;
wire _00848_;
wire _00849_;
wire _00850_;
wire _00851_;
wire _00852_;
wire _00853_;
wire _00854_;
wire _00855_;
wire _00856_;
wire _00857_;
wire _00858_;
wire _00859_;
wire _00860_;
wire _00861_;
wire _00862_;
wire _00863_;
wire _00864_;
wire _00865_;
wire _00866_;
wire _00867_;
wire _00868_;
wire _00869_;
wire _00870_;
wire _00871_;
wire _00872_;
wire _00873_;
wire _00874_;
wire _00875_;
wire _00876_;
wire _00877_;
wire _00878_;
wire _00879_;
wire _00880_;
wire _00881_;
wire _00882_;
wire _00883_;
wire _00884_;
wire _00885_;
wire _00886_;
wire _00887_;
wire _00888_;
wire _00889_;
wire _00890_;
wire _00891_;
wire _00892_;
wire _00893_;
wire _00894_;
wire _00895_;
wire _00896_;
wire _00897_;
wire _00898_;
wire _00899_;
wire _00900_;
wire _00901_;
wire _00902_;
wire _00903_;
wire _00904_;
wire _00905_;
wire _00906_;
wire _00907_;
wire _00908_;
wire _00909_;
wire _00910_;
wire _00911_;
wire _00912_;
wire _00913_;
wire _00914_;
wire _00915_;
wire _00916_;
wire _00917_;
wire _00918_;
wire _00919_;
wire _00920_;
wire _00921_;
wire _00922_;
wire _00923_;
wire _00924_;
wire _00925_;
wire _00926_;
wire _00927_;
wire _00928_;
wire _00929_;
wire _00930_;
wire _00931_;
wire _00932_;
wire _00933_;
wire _00934_;
wire _00935_;
wire _00936_;
wire _00937_;
wire _00938_;
wire _00939_;
wire _00940_;
wire _00941_;
wire _00942_;
wire _00943_;
wire _00944_;
wire _00945_;
wire _00946_;
wire _00947_;
wire _00948_;
wire _00949_;
wire _00950_;
wire _00951_;
wire _00952_;
wire _00953_;
wire _00954_;
wire _00955_;
wire _00956_;
wire _00957_;
wire _00958_;
wire _00959_;
wire _00960_;
wire _00961_;
wire _00962_;
wire _00963_;
wire _00964_;
wire _00965_;
wire _00966_;
wire _00967_;
wire _00968_;
wire _00969_;
wire _00970_;
wire _00971_;
wire _00972_;
wire _00973_;
wire _00974_;
wire _00975_;
wire _00976_;
wire _00977_;
wire _00978_;
wire _00979_;
wire _00980_;
wire _00981_;
wire _00982_;
wire _00983_;
wire _00984_;
wire _00985_;
wire _00986_;
wire _00987_;
wire _00988_;
wire _00989_;
wire _00990_;
wire _00991_;
wire _00992_;
wire _00993_;
wire _00994_;
wire _00995_;
wire _00996_;
wire _00997_;
wire _00998_;
wire _00999_;
wire _01000_;
wire _01001_;
wire _01002_;
wire _01003_;
wire _01004_;
wire _01005_;
wire _01006_;
wire _01007_;
wire _01008_;
wire _01009_;
wire _01010_;
wire _01011_;
wire _01012_;
wire _01013_;
wire _01014_;
wire _01015_;
wire _01016_;
wire _01017_;
wire _01018_;
wire _01019_;
wire _01020_;
wire _01021_;
wire _01022_;
wire _01023_;
wire _01024_;
wire _01025_;
wire _01026_;
wire _01027_;
wire _01028_;
wire _01029_;
wire _01030_;
wire _01031_;
wire _01032_;
wire _01033_;
wire _01034_;
wire _01035_;
wire _01036_;
wire _01037_;
wire _01038_;
wire _01039_;
wire _01040_;
wire _01041_;
wire _01042_;
wire _01043_;
wire _01044_;
wire _01045_;
wire _01046_;
wire _01047_;
wire _01048_;
wire _01049_;
wire _01050_;
wire _01051_;
wire _01052_;
wire _01053_;
wire _01054_;
wire _01055_;
wire _01056_;
wire _01057_;
wire _01058_;
wire _01059_;
wire _01060_;
wire _01061_;
wire _01062_;
wire _01063_;
wire _01064_;
wire _01065_;
wire _01066_;
wire _01067_;
wire _01068_;
wire _01069_;
wire _01070_;
wire _01071_;
wire _01072_;
wire _01073_;
wire _01074_;
wire _01075_;
wire _01076_;
wire _01077_;
wire _01078_;
wire _01079_;
wire _01080_;
wire _01081_;
wire _01082_;
wire _01083_;
wire _01084_;
wire _01085_;
wire _01086_;
wire _01087_;
wire _01088_;
wire _01089_;
wire _01090_;
wire _01091_;
wire _01092_;
wire _01093_;
wire _01094_;
wire _01095_;
wire _01096_;
wire _01097_;
wire _01098_;
wire _01099_;
wire _01100_;
wire _01101_;
wire _01102_;
wire _01103_;
wire _01104_;
wire _01105_;
wire _01106_;
wire _01107_;
wire _01108_;
wire _01109_;
wire _01110_;
wire _01111_;
wire _01112_;
wire _01113_;
wire _01114_;
wire _01115_;
wire _01116_;
wire _01117_;
wire _01118_;
wire _01119_;
wire _01120_;
wire _01121_;
wire _01122_;
wire _01123_;
wire _01124_;
wire _01125_;
wire _01126_;
wire _01127_;
wire _01128_;
wire _01129_;
wire _01130_;
wire _01131_;
wire _01132_;
wire _01133_;
wire _01134_;
wire _01135_;
wire _01136_;
wire _01137_;
wire _01138_;
wire _01139_;
wire _01140_;
wire _01141_;
wire _01142_;
wire _01143_;
wire _01144_;
wire _01145_;
wire _01146_;
wire _01147_;
wire _01148_;
wire _01149_;
wire _01150_;
wire _01151_;
wire _01152_;
wire _01153_;
wire _01154_;
wire _01155_;
wire _01156_;
wire _01157_;
wire _01158_;
wire _01159_;
wire _01160_;
wire _01161_;
wire _01162_;
wire _01163_;
wire _01164_;
wire _01165_;
wire _01166_;
wire _01167_;
wire _01168_;
wire _01169_;
wire _01170_;
wire _01171_;
wire _01172_;
wire _01173_;
wire _01174_;
wire _01175_;
wire _01176_;
wire _01177_;
wire _01178_;
wire _01179_;
wire _01180_;
wire _01181_;
wire _01182_;
wire _01183_;
wire _01184_;
wire _01185_;
wire _01186_;
wire _01187_;
wire _01188_;
wire _01189_;
wire _01190_;
wire _01191_;
wire _01192_;
wire _01193_;
wire _01194_;
wire _01195_;
wire _01196_;
wire _01197_;
wire _01198_;
wire _01199_;
wire _01200_;
wire _01201_;
wire _01202_;
wire _01203_;
wire _01204_;
wire _01205_;
wire _01206_;
wire _01207_;
wire _01208_;
wire _01209_;
wire _01210_;
wire _01211_;
wire _01212_;
wire _01213_;
wire _01214_;
wire _01215_;
wire _01216_;
wire _01217_;
wire _01218_;
wire _01219_;
wire _01220_;
wire _01221_;
wire _01222_;
wire _01223_;
wire _01224_;
wire _01225_;
wire _01226_;
wire _01227_;
wire _01228_;
wire _01229_;
wire _01230_;
wire _01231_;
wire _01232_;
wire _01233_;
wire _01234_;
wire _01235_;
wire _01236_;
wire _01237_;
wire _01238_;
wire _01239_;
wire _01240_;
wire _01241_;
wire _01242_;
wire _01243_;
wire _01244_;
wire _01245_;
wire _01246_;
wire _01247_;
wire _01248_;
wire _01249_;
wire _01250_;
wire _01251_;
wire _01252_;
wire _01253_;
wire _01254_;
wire _01255_;
wire _01256_;
wire _01257_;
wire _01258_;
wire _01259_;
wire _01260_;
wire _01261_;
wire _01262_;
wire _01263_;
wire _01264_;
wire _01265_;
wire _01266_;
wire _01267_;
wire _01268_;
wire _01269_;
wire _01270_;
wire _01271_;
wire _01272_;
wire _01273_;
wire _01274_;
wire _01275_;
wire _01276_;
wire _01277_;
wire _01278_;
wire _01279_;
wire _01280_;
wire _01281_;
wire _01282_;
wire _01283_;
wire _01284_;
wire _01285_;
wire _01286_;
wire _01287_;
wire _01288_;
wire _01289_;
wire _01290_;
wire _01291_;
wire _01292_;
wire _01293_;
wire _01294_;
wire _01295_;
wire _01296_;
wire _01297_;
wire _01298_;
wire _01299_;
wire _01300_;
wire _01301_;
wire _01302_;
wire _01303_;
wire _01304_;
wire _01305_;
wire _01306_;
wire _01307_;
wire _01308_;
wire _01309_;
wire _01310_;
wire _01311_;
wire _01312_;
wire _01313_;
wire _01314_;
wire _01315_;
wire _01316_;
wire _01317_;
wire _01318_;
wire _01319_;
wire _01320_;
wire _01321_;
wire _01322_;
wire _01323_;
wire _01324_;
wire _01325_;
wire _01326_;
wire _01327_;
wire _01328_;
wire _01329_;
wire _01330_;
wire _01331_;
wire _01332_;
wire _01333_;
wire _01334_;
wire _01335_;
wire _01336_;
wire _01337_;
wire _01338_;
wire _01339_;
wire _01340_;
wire _01341_;
wire _01342_;
wire _01343_;
wire _01344_;
wire _01345_;
wire _01346_;
wire _01347_;
wire _01348_;
wire _01349_;
wire _01350_;
wire _01351_;
wire _01352_;
wire _01353_;
wire _01354_;
wire _01355_;
wire _01356_;
wire _01357_;
wire _01358_;
wire _01359_;
wire _01360_;
wire _01361_;
wire _01362_;
wire _01363_;
wire _01364_;
wire _01365_;
wire _01366_;
wire _01367_;
wire _01368_;
wire _01369_;
wire _01370_;
wire _01371_;
wire _01372_;
wire _01373_;
wire _01374_;
wire _01375_;
wire _01376_;
wire _01377_;
wire _01378_;
wire _01379_;
wire _01380_;
wire _01381_;
wire _01382_;
wire _01383_;
wire _01384_;
wire _01385_;
wire _01386_;
wire _01387_;
wire _01388_;
wire _01389_;
wire _01390_;
wire _01391_;
wire _01392_;
wire _01393_;
wire _01394_;
wire _01395_;
wire _01396_;
wire _01397_;
wire _01398_;
wire _01399_;
wire _01400_;
wire _01401_;
wire _01402_;
wire _01403_;
wire _01404_;
wire _01405_;
wire _01406_;
wire _01407_;
wire _01408_;
wire _01409_;
wire _01410_;
wire _01411_;
wire _01412_;
wire _01413_;
wire _01414_;
wire _01415_;
wire _01416_;
wire _01417_;
wire _01418_;
wire _01419_;
wire _01420_;
wire _01421_;
wire _01422_;
wire _01423_;
wire _01424_;
wire _01425_;
wire _01426_;
wire _01427_;
wire _01428_;
wire _01429_;
wire _01430_;
wire _01431_;
wire _01432_;
wire _01433_;
wire _01434_;
wire _01435_;
wire _01436_;
wire _01437_;
wire _01438_;
wire _01439_;
wire _01440_;
wire _01441_;
wire _01442_;
wire _01443_;
wire _01444_;
wire _01445_;
wire _01446_;
wire _01447_;
wire _01448_;
wire _01449_;
wire _01450_;
wire _01451_;
wire _01452_;
wire _01453_;
wire _01454_;
wire _01455_;
wire _01456_;
wire _01457_;
wire _01458_;
wire _01459_;
wire _01460_;
wire _01461_;
wire _01462_;
wire _01463_;
wire _01464_;
wire _01465_;
wire _01466_;
wire _01467_;
wire _01468_;
wire _01469_;
wire _01470_;
wire _01471_;
wire _01472_;
wire _01473_;
wire _01474_;
wire _01475_;
wire _01476_;
wire _01477_;
wire _01478_;
wire _01479_;
wire _01480_;
wire _01481_;
wire _01482_;
wire _01483_;
wire _01484_;
wire _01485_;
wire _01486_;
wire _01487_;
wire _01488_;
wire _01489_;
wire _01490_;
wire _01491_;
wire _01492_;
wire _01493_;
wire _01494_;
wire _01495_;
wire _01496_;
wire _01497_;
wire _01498_;
wire _01499_;
wire _01500_;
wire _01501_;
wire _01502_;
wire _01503_;
wire _01504_;
wire _01505_;
wire _01506_;
wire _01507_;
wire _01508_;
wire _01509_;
wire _01510_;
wire _01511_;
wire _01512_;
wire _01513_;
wire _01514_;
wire _01515_;
wire _01516_;
wire _01517_;
wire _01518_;
wire _01519_;
wire _01520_;
wire _01521_;
wire _01522_;
wire _01523_;
wire _01524_;
wire _01525_;
wire _01526_;
wire _01527_;
wire _01528_;
wire _01529_;
wire _01530_;
wire _01531_;
wire _01532_;
wire _01533_;
wire _01534_;
wire _01535_;
wire _01536_;
wire _01537_;
wire _01538_;
wire _01539_;
wire _01540_;
wire _01541_;
wire _01542_;
wire _01543_;
wire _01544_;
wire _01545_;
wire _01546_;
wire _01547_;
wire _01548_;
wire _01549_;
wire _01550_;
wire _01551_;
wire _01552_;
wire _01553_;
wire _01554_;
wire _01555_;
wire _01556_;
wire _01557_;
wire _01558_;
wire _01559_;
wire _01560_;
wire _01561_;
wire _01562_;
wire _01563_;
wire _01564_;
wire _01565_;
wire _01566_;
wire _01567_;
wire _01568_;
wire _01569_;
wire _01570_;
wire _01571_;
wire _01572_;
wire _01573_;
wire _01574_;
wire _01575_;
wire _01576_;
wire _01577_;
wire _01578_;
wire _01579_;
wire _01580_;
wire _01581_;
wire _01582_;
wire _01583_;
wire _01584_;
wire _01585_;
wire _01586_;
wire _01587_;
wire _01588_;
wire _01589_;
wire _01590_;
wire _01591_;
wire _01592_;
wire _01593_;
wire _01594_;
wire _01595_;
wire _01596_;
wire _01597_;
wire _01598_;
wire _01599_;
wire _01600_;
wire _01601_;
wire _01602_;
wire _01603_;
wire _01604_;
wire _01605_;
wire _01606_;
wire _01607_;
wire _01608_;
wire _01609_;
wire _01610_;
wire _01611_;
wire _01612_;
wire _01613_;
wire _01614_;
wire _01615_;
wire _01616_;
wire _01617_;
wire _01618_;
wire _01619_;
wire _01620_;
wire _01621_;
wire _01622_;
wire _01623_;
wire _01624_;
wire _01625_;
wire _01626_;
wire _01627_;
wire _01628_;
wire _01629_;
wire _01630_;
wire _01631_;
wire _01632_;
wire _01633_;
wire _01634_;
wire _01635_;
wire _01636_;
wire _01637_;
wire _01638_;
wire _01639_;
wire _01640_;
wire _01641_;
wire _01642_;
wire _01643_;
wire _01644_;
wire _01645_;
wire _01646_;
wire _01647_;
wire _01648_;
wire _01649_;
wire _01650_;
wire _01651_;
wire _01652_;
wire _01653_;
wire _01654_;
wire _01655_;
wire _01656_;
wire _01657_;
wire _01658_;
wire _01659_;
wire _01660_;
wire _01661_;
wire _01662_;
wire _01663_;
wire _01664_;
wire _01665_;
wire _01666_;
wire _01667_;
wire _01668_;
wire _01669_;
wire _01670_;
wire _01671_;
wire _01672_;
wire _01673_;
wire _01674_;
wire _01675_;
wire _01676_;
wire _01677_;
wire _01678_;
wire _01679_;
wire _01680_;
wire _01681_;
wire _01682_;
wire _01683_;
wire _01684_;
wire _01685_;
wire _01686_;
wire _01687_;
wire _01688_;
wire _01689_;
wire _01690_;
wire _01691_;
wire _01692_;
wire _01693_;
wire _01694_;
wire _01695_;
wire _01696_;
wire _01697_;
wire _01698_;
wire _01699_;
wire _01700_;
wire _01701_;
wire _01702_;
wire _01703_;
wire _01704_;
wire _01705_;
wire _01706_;
wire _01707_;
wire _01708_;
wire _01709_;
wire _01710_;
wire _01711_;
wire _01712_;
wire _01713_;
wire _01714_;
wire _01715_;
wire _01716_;
wire _01717_;
wire _01718_;
wire _01719_;
wire _01720_;
wire _01721_;
wire _01722_;
wire _01723_;
wire _01724_;
wire _01725_;
wire _01726_;
wire _01727_;
wire _01728_;
wire _01729_;
wire _01730_;
wire _01731_;
wire _01732_;
wire _01733_;
wire _01734_;
wire _01735_;
wire _01736_;
wire _01737_;
wire _01738_;
wire _01739_;
wire _01740_;
wire _01741_;
wire _01742_;
wire _01743_;
wire _01744_;
wire _01745_;
wire _01746_;
wire _01747_;
wire _01748_;
wire _01749_;
wire _01750_;
wire _01751_;
wire _01752_;
wire _01753_;
wire _01754_;
wire _01755_;
wire _01756_;
wire _01757_;
wire _01758_;
wire _01759_;
wire _01760_;
wire _01761_;
wire _01762_;
wire _01763_;
wire _01764_;
wire _01765_;
wire _01766_;
wire _01767_;
wire _01768_;
wire _01769_;
wire _01770_;
wire _01771_;
wire _01772_;
wire _01773_;
wire _01774_;
wire _01775_;
wire _01776_;
wire _01777_;
wire _01778_;
wire _01779_;
wire _01780_;
wire _01781_;
wire _01782_;
wire _01783_;
wire _01784_;
wire _01785_;
wire _01786_;
wire _01787_;
wire _01788_;
wire _01789_;
wire _01790_;
wire _01791_;
wire _01792_;
wire _01793_;
wire _01794_;
wire _01795_;
wire _01796_;
wire _01797_;
wire _01798_;
wire _01799_;
wire _01800_;
wire _01801_;
wire _01802_;
wire _01803_;
wire _01804_;
wire _01805_;
wire _01806_;
wire _01807_;
wire _01808_;
wire _01809_;
wire _01810_;
wire _01811_;
wire _01812_;
wire _01813_;
wire _01814_;
wire _01815_;
wire _01816_;
wire _01817_;
wire _01818_;
wire _01819_;
wire _01820_;
wire _01821_;
wire _01822_;
wire _01823_;
wire _01824_;
wire _01825_;
wire _01826_;
wire _01827_;
wire _01828_;
wire _01829_;
wire _01830_;
wire _01831_;
wire _01832_;
wire _01833_;
wire _01834_;
wire _01835_;
wire _01836_;
wire _01837_;
wire _01838_;
wire _01839_;
wire _01840_;
wire _01841_;
wire _01842_;
wire _01843_;
wire _01844_;
wire _01845_;
wire _01846_;
wire _01847_;
wire _01848_;
wire _01849_;
wire _01850_;
wire _01851_;
wire _01852_;
wire _01853_;
wire _01854_;
wire _01855_;
wire _01856_;
wire _01857_;
wire _01858_;
wire _01859_;
wire _01860_;
wire _01861_;
wire _01862_;
wire _01863_;
wire _01864_;
wire _01865_;
wire _01866_;
wire _01867_;
wire _01868_;
wire _01869_;
wire _01870_;
wire _01871_;
wire _01872_;
wire _01873_;
wire _01874_;
wire _01875_;
wire _01876_;
wire _01877_;
wire _01878_;
wire _01879_;
wire _01880_;
wire _01881_;
wire _01882_;
wire _01883_;
wire _01884_;
wire _01885_;
wire _01886_;
wire _01887_;
wire _01888_;
wire _01889_;
wire _01890_;
wire _01891_;
wire _01892_;
wire _01893_;
wire _01894_;
wire _01895_;
wire _01896_;
wire _01897_;
wire _01898_;
wire _01899_;
wire _01900_;
wire _01901_;
wire _01902_;
wire _01903_;
wire _01904_;
wire _01905_;
wire _01906_;
wire _01907_;
wire _01908_;
wire _01909_;
wire _01910_;
wire _01911_;
wire _01912_;
wire _01913_;
wire _01914_;
wire _01915_;
wire _01916_;
wire _01917_;
wire _01918_;
wire _01919_;
wire _01920_;
wire _01921_;
wire _01922_;
wire _01923_;
wire _01924_;
wire _01925_;
wire _01926_;
wire _01927_;
wire _01928_;
wire _01929_;
wire _01930_;
wire _01931_;
wire _01932_;
wire _01933_;
wire _01934_;
wire _01935_;
wire _01936_;
wire _01937_;
wire _01938_;
wire _01939_;
wire _01940_;
wire _01941_;
wire _01942_;
wire _01943_;
wire _01944_;
wire _01945_;
wire _01946_;
wire _01947_;
wire _01948_;
wire _01949_;
wire _01950_;
wire _01951_;
wire _01952_;
wire _01953_;
wire _01954_;
wire _01955_;
wire _01956_;
wire _01957_;
wire _01958_;
wire _01959_;
wire _01960_;
wire _01961_;
wire _01962_;
wire _01963_;
wire _01964_;
wire _01965_;
wire _01966_;
wire _01967_;
wire _01968_;
wire _01969_;
wire _01970_;
wire _01971_;
wire _01972_;
wire _01973_;
wire _01974_;
wire _01975_;
wire _01976_;
wire _01977_;
wire _01978_;
wire _01979_;
wire _01980_;
wire _01981_;
wire _01982_;
wire _01983_;
wire _01984_;
wire _01985_;
wire _01986_;
wire _01987_;
wire _01988_;
wire _01989_;
wire _01990_;
wire _01991_;
wire _01992_;
wire _01993_;
wire _01994_;
wire _01995_;
wire _01996_;
wire _01997_;
wire _01998_;
wire _01999_;
wire _02000_;
wire _02001_;
wire _02002_;
wire _02003_;
wire _02004_;
wire _02005_;
wire _02006_;
wire _02007_;
wire _02008_;
wire _02009_;
wire _02010_;
wire _02011_;
wire _02012_;
wire _02013_;
wire _02014_;
wire _02015_;
wire _02016_;
wire _02017_;
wire _02018_;
wire _02019_;
wire _02020_;
wire _02021_;
wire _02022_;
wire _02023_;
wire _02024_;
wire _02025_;
wire _02026_;
wire _02027_;
wire _02028_;
wire _02029_;
wire _02030_;
wire _02031_;
wire _02032_;
wire _02033_;
wire _02034_;
wire _02035_;
wire _02036_;
wire _02037_;
wire _02038_;
wire _02039_;
wire _02040_;
wire _02041_;
wire _02042_;
wire _02043_;
wire _02044_;
wire _02045_;
wire _02046_;
wire _02047_;
wire _02048_;
wire _02049_;
wire _02050_;
wire _02051_;
wire _02052_;
wire _02053_;
wire _02054_;
wire _02055_;
wire _02056_;
wire _02057_;
wire _02058_;
wire _02059_;
wire _02060_;
wire _02061_;
wire _02062_;
wire _02063_;
wire _02064_;
wire _02065_;
wire _02066_;
wire _02067_;
wire _02068_;
wire _02069_;
wire _02070_;
wire _02071_;
wire _02072_;
wire _02073_;
wire _02074_;
wire _02075_;
wire _02076_;
wire _02077_;
wire _02078_;
wire _02079_;
wire _02080_;
wire _02081_;
wire _02082_;
wire _02083_;
wire _02084_;
wire _02085_;
wire _02086_;
wire _02087_;
wire _02088_;
wire _02089_;
wire _02090_;
wire _02091_;
wire _02092_;
wire _02093_;
wire _02094_;
wire _02095_;
wire _02096_;
wire _02097_;
wire _02098_;
wire _02099_;
wire _02100_;
wire _02101_;
wire _02102_;
wire _02103_;
wire _02104_;
wire _02105_;
wire _02106_;
wire _02107_;
wire _02108_;
wire _02109_;
wire _02110_;
wire _02111_;
wire _02112_;
wire _02113_;
wire _02114_;
wire _02115_;
wire _02116_;
wire _02117_;
wire _02118_;
wire _02119_;
wire _02120_;
wire _02121_;
wire _02122_;
wire _02123_;
wire _02124_;
wire _02125_;
wire _02126_;
wire _02127_;
wire _02128_;
wire _02129_;
wire _02130_;
wire _02131_;
wire _02132_;
wire _02133_;
wire _02134_;
wire _02135_;
wire _02136_;
wire _02137_;
wire _02138_;
wire _02139_;
wire _02140_;
wire _02141_;
wire _02142_;
wire _02143_;
wire _02144_;
wire _02145_;
wire _02146_;
wire _02147_;
wire _02148_;
wire _02149_;
wire _02150_;
wire _02151_;
wire _02152_;
wire _02153_;
wire _02154_;
wire _02155_;
wire _02156_;
wire _02157_;
wire _02158_;
wire _02159_;
wire _02160_;
wire _02161_;
wire _02162_;
wire _02163_;
wire _02164_;
wire _02165_;
wire _02166_;
wire _02167_;
wire _02168_;
wire _02169_;
wire _02170_;
wire _02171_;
wire _02172_;
wire _02173_;
wire _02174_;
wire _02175_;
wire _02176_;
wire _02177_;
wire _02178_;
wire _02179_;
wire _02180_;
wire _02181_;
wire _02182_;
wire _02183_;
wire _02184_;
wire _02185_;
wire _02186_;
wire _02187_;
wire _02188_;
wire _02189_;
wire _02190_;
wire _02191_;
wire _02192_;
wire _02193_;
wire _02194_;
wire _02195_;
wire _02196_;
wire _02197_;
wire _02198_;
wire _02199_;
wire _02200_;
wire _02201_;
wire _02202_;
wire _02203_;
wire _02204_;
wire _02205_;
wire _02206_;
wire _02207_;
wire _02208_;
wire _02209_;
wire _02210_;
wire _02211_;
wire _02212_;
wire _02213_;
wire _02214_;
wire _02215_;
wire _02216_;
wire _02217_;
wire _02218_;
wire _02219_;
wire _02220_;
wire _02221_;
wire _02222_;
wire _02223_;
wire _02224_;
wire _02225_;
wire _02226_;
wire _02227_;
wire _02228_;
wire _02229_;
wire _02230_;
wire _02231_;
wire _02232_;
wire _02233_;
wire _02234_;
wire _02235_;
wire _02236_;
wire _02237_;
wire _02238_;
wire _02239_;
wire _02240_;
wire _02241_;
wire _02242_;
wire _02243_;
wire _02244_;
wire _02245_;
wire _02246_;
wire _02247_;
wire _02248_;
wire _02249_;
wire _02250_;
wire _02251_;
wire _02252_;
wire _02253_;
wire _02254_;
wire _02255_;
wire _02256_;
wire _02257_;
wire _02258_;
wire _02259_;
wire _02260_;
wire _02261_;
wire _02262_;
wire _02263_;
wire _02264_;
wire _02265_;
wire _02266_;
wire _02267_;
wire _02268_;
wire _02269_;
wire _02270_;
wire _02271_;
wire _02272_;
wire _02273_;
wire _02274_;
wire _02275_;
wire _02276_;
wire _02277_;
wire _02278_;
wire _02279_;
wire _02280_;
wire _02281_;
wire _02282_;
wire _02283_;
wire _02284_;
wire _02285_;
wire _02286_;
wire _02287_;
wire _02288_;
wire _02289_;
wire _02290_;
wire _02291_;
wire _02292_;
wire _02293_;
wire _02294_;
wire _02295_;
wire _02296_;
wire _02297_;
wire _02298_;
wire _02299_;
wire _02300_;
wire _02301_;
wire _02302_;
wire _02303_;
wire _02304_;
wire _02305_;
wire _02306_;
wire _02307_;
wire _02308_;
wire _02309_;
wire _02310_;
wire _02311_;
wire _02312_;
wire _02313_;
wire _02314_;
wire _02315_;
wire _02316_;
wire _02317_;
wire _02318_;
wire _02319_;
wire _02320_;
wire _02321_;
wire _02322_;
wire _02323_;
wire _02324_;
wire _02325_;
wire _02326_;
wire _02327_;
wire _02328_;
wire _02329_;
wire _02330_;
wire _02331_;
wire _02332_;
wire _02333_;
wire _02334_;
wire _02335_;
wire _02336_;
wire _02337_;
wire _02338_;
wire _02339_;
wire _02340_;
wire _02341_;
wire _02342_;
wire _02343_;
wire _02344_;
wire _02345_;
wire _02346_;
wire _02347_;
wire _02348_;
wire _02349_;
wire _02350_;
wire _02351_;
wire _02352_;
wire _02353_;
wire _02354_;
wire _02355_;
wire _02356_;
wire _02357_;
wire _02358_;
wire _02359_;
wire _02360_;
wire _02361_;
wire _02362_;
wire _02363_;
wire _02364_;
wire _02365_;
wire _02366_;
wire _02367_;
wire _02368_;
wire _02369_;
wire _02370_;
wire _02371_;
wire _02372_;
wire _02373_;
wire _02374_;
wire _02375_;
wire _02376_;
wire _02377_;
wire _02378_;
wire _02379_;
wire _02380_;
wire _02381_;
wire _02382_;
wire _02383_;
wire _02384_;
wire _02385_;
wire _02386_;
wire _02387_;
wire _02388_;
wire _02389_;
wire _02390_;
wire _02391_;
wire _02392_;
wire _02393_;
wire _02394_;
wire _02395_;
wire _02396_;
wire _02397_;
wire _02398_;
wire _02399_;
wire _02400_;
wire _02401_;
wire _02402_;
wire _02403_;
wire _02404_;
wire _02405_;
wire _02406_;
wire _02407_;
wire _02408_;
wire _02409_;
wire _02410_;
wire _02411_;
wire _02412_;
wire _02413_;
wire _02414_;
wire _02415_;
wire _02416_;
wire _02417_;
wire _02418_;
wire _02419_;
wire _02420_;
wire _02421_;
wire _02422_;
wire _02423_;
wire _02424_;
wire _02425_;
wire _02426_;
wire _02427_;
wire _02428_;
wire _02429_;
wire _02430_;
wire _02431_;
wire _02432_;
wire _02433_;
wire _02434_;
wire _02435_;
wire _02436_;
wire _02437_;
wire _02438_;
wire _02439_;
wire _02440_;
wire _02441_;
wire _02442_;
wire _02443_;
wire _02444_;
wire _02445_;
wire _02446_;
wire _02447_;
wire _02448_;
wire _02449_;
wire _02450_;
wire _02451_;
wire _02452_;
wire _02453_;
wire _02454_;
wire _02455_;
wire _02456_;
wire _02457_;
wire _02458_;
wire _02459_;
wire _02460_;
wire _02461_;
wire _02462_;
wire _02463_;
wire _02464_;
wire _02465_;
wire _02466_;
wire _02467_;
wire _02468_;
wire _02469_;
wire _02470_;
wire _02471_;
wire _02472_;
wire _02473_;
wire _02474_;
wire _02475_;
wire _02476_;
wire _02477_;
wire _02478_;
wire _02479_;
wire _02480_;
wire _02481_;
wire _02482_;
wire _02483_;
wire _02484_;
wire _02485_;
wire _02486_;
wire _02487_;
wire _02488_;
wire _02489_;
wire _02490_;
wire _02491_;
wire _02492_;
wire _02493_;
wire _02494_;
wire _02495_;
wire _02496_;
wire _02497_;
wire _02498_;
wire _02499_;
wire _02500_;
wire _02501_;
wire _02502_;
wire _02503_;
wire _02504_;
wire _02505_;
wire _02506_;
wire _02507_;
wire _02508_;
wire _02509_;
wire _02510_;
wire _02511_;
wire _02512_;
wire _02513_;
wire _02514_;
wire _02515_;
wire _02516_;
wire _02517_;
wire _02518_;
wire _02519_;
wire _02520_;
wire _02521_;
wire _02522_;
wire _02523_;
wire _02524_;
wire _02525_;
wire _02526_;
wire _02527_;
wire _02528_;
wire _02529_;
wire _02530_;
wire _02531_;
wire _02532_;
wire _02533_;
wire _02534_;
wire _02535_;
wire _02536_;
wire _02537_;
wire _02538_;
wire _02539_;
wire _02540_;
wire _02541_;
wire _02542_;
wire _02543_;
wire _02544_;
wire _02545_;
wire _02546_;
wire _02547_;
wire _02548_;
wire _02549_;
wire _02550_;
wire _02551_;
wire _02552_;
wire _02553_;
wire _02554_;
wire _02555_;
wire _02556_;
wire _02557_;
wire _02558_;
wire _02559_;
wire _02560_;
wire _02561_;
wire _02562_;
wire _02563_;
wire _02564_;
wire _02565_;
wire _02566_;
wire _02567_;
wire _02568_;
wire _02569_;
wire _02570_;
wire _02571_;
wire _02572_;
wire _02573_;
wire _02574_;
wire _02575_;
wire _02576_;
wire _02577_;
wire _02578_;
wire _02579_;
wire _02580_;
wire _02581_;
wire _02582_;
wire _02583_;
wire _02584_;
wire _02585_;
wire _02586_;
wire _02587_;
wire _02588_;
wire _02589_;
wire _02590_;
wire _02591_;
wire _02592_;
wire _02593_;
wire _02594_;
wire _02595_;
wire _02596_;
wire _02597_;
wire _02598_;
wire _02599_;
wire _02600_;
wire _02601_;
wire _02602_;
wire _02603_;
wire _02604_;
wire _02605_;
wire _02606_;
wire _02607_;
wire _02608_;
wire _02609_;
wire _02610_;
wire _02611_;
wire _02612_;
wire _02613_;
wire _02614_;
wire _02615_;
wire _02616_;
wire _02617_;
wire _02618_;
wire _02619_;
wire _02620_;
wire _02621_;
wire _02622_;
wire _02623_;
wire _02624_;
wire _02625_;
wire _02626_;
wire _02627_;
wire _02628_;
wire _02629_;
wire _02630_;
wire _02631_;
wire _02632_;
wire _02633_;
wire _02634_;
wire _02635_;
wire _02636_;
wire _02637_;
wire _02638_;
wire _02639_;
wire _02640_;
wire _02641_;
wire _02642_;
wire _02643_;
wire _02644_;
wire _02645_;
wire _02646_;
wire _02647_;
wire _02648_;
wire _02649_;
wire _02650_;
wire _02651_;
wire _02652_;
wire _02653_;
wire _02654_;
wire _02655_;
wire _02656_;
wire _02657_;
wire _02658_;
wire _02659_;
wire _02660_;
wire _02661_;
wire _02662_;
wire _02663_;
wire _02664_;
wire _02665_;
wire _02666_;
wire _02667_;
wire _02668_;
wire _02669_;
wire _02670_;
wire _02671_;
wire _02672_;
wire _02673_;
wire _02674_;
wire _02675_;
wire _02676_;
wire _02677_;
wire _02678_;
wire _02679_;
wire _02680_;
wire _02681_;
wire _02682_;
wire _02683_;
wire _02684_;
wire _02685_;
wire _02686_;
wire _02687_;
wire _02688_;
wire _02689_;
wire _02690_;
wire _02691_;
wire _02692_;
wire _02693_;
wire _02694_;
wire _02695_;
wire _02696_;
wire _02697_;
wire _02698_;
wire _02699_;
wire _02700_;
wire _02701_;
wire _02702_;
wire _02703_;
wire _02704_;
wire _02705_;
wire _02706_;
wire _02707_;
wire _02708_;
wire _02709_;
wire _02710_;
wire _02711_;
wire _02712_;
wire _02713_;
wire _02714_;
wire _02715_;
wire _02716_;
wire _02717_;
wire _02718_;
wire _02719_;
wire _02720_;
wire _02721_;
wire _02722_;
wire _02723_;
wire _02724_;
wire _02725_;
wire _02726_;
wire _02727_;
wire _02728_;
wire _02729_;
wire _02730_;
wire _02731_;
wire _02732_;
wire _02733_;
wire _02734_;
wire _02735_;
wire _02736_;
wire _02737_;
wire _02738_;
wire _02739_;
wire _02740_;
wire _02741_;
wire _02742_;
wire _02743_;
wire _02744_;
wire _02745_;
wire _02746_;
wire _02747_;
wire _02748_;
wire _02749_;
wire _02750_;
wire _02751_;
wire _02752_;
wire _02753_;
wire _02754_;
wire _02755_;
wire _02756_;
wire _02757_;
wire _02758_;
wire _02759_;
wire _02760_;
wire _02761_;
wire _02762_;
wire _02763_;
wire _02764_;
wire _02765_;
wire _02766_;
wire _02767_;
wire _02768_;
wire _02769_;
wire _02770_;
wire _02771_;
wire _02772_;
wire _02773_;
wire _02774_;
wire _02775_;
wire _02776_;
wire _02777_;
wire _02778_;
wire _02779_;
wire _02780_;
wire _02781_;
wire _02782_;
wire _02783_;
wire _02784_;
wire _02785_;
wire _02786_;
wire _02787_;
wire _02788_;
wire _02789_;
wire _02790_;
wire _02791_;
wire _02792_;
wire _02793_;
wire _02794_;
wire _02795_;
wire _02796_;
wire _02797_;
wire _02798_;
wire _02799_;
wire _02800_;
wire _02801_;
wire _02802_;
wire _02803_;
wire _02804_;
wire _02805_;
wire _02806_;
wire _02807_;
wire _02808_;
wire _02809_;
wire _02810_;
wire _02811_;
wire _02812_;
wire _02813_;
wire _02814_;
wire _02815_;
wire _02816_;
wire _02817_;
wire _02818_;
wire _02819_;
wire _02820_;
wire _02821_;
wire _02822_;
wire _02823_;
wire _02824_;
wire _02825_;
wire _02826_;
wire _02827_;
wire _02828_;
wire _02829_;
wire _02830_;
wire _02831_;
wire _02832_;
wire _02833_;
wire _02834_;
wire _02835_;
wire _02836_;
wire _02837_;
wire _02838_;
wire _02839_;
wire _02840_;
wire _02841_;
wire _02842_;
wire _02843_;
wire _02844_;
wire _02845_;
wire _02846_;
wire _02847_;
wire _02848_;
wire _02849_;
wire _02850_;
wire _02851_;
wire _02852_;
wire _02853_;
wire _02854_;
wire _02855_;
wire _02856_;
wire _02857_;
wire _02858_;
wire _02859_;
wire _02860_;
wire _02861_;
wire _02862_;
wire _02863_;
wire _02864_;
wire _02865_;
wire _02866_;
wire _02867_;
wire _02868_;
wire _02869_;
wire _02870_;
wire _02871_;
wire _02872_;
wire _02873_;
wire _02874_;
wire _02875_;
wire _02876_;
wire _02877_;
wire _02878_;
wire _02879_;
wire _02880_;
wire _02881_;
wire _02882_;
wire _02883_;
wire _02884_;
wire _02885_;
wire _02886_;
wire _02887_;
wire _02888_;
wire _02889_;
wire _02890_;
wire _02891_;
wire _02892_;
wire _02893_;
wire _02894_;
wire _02895_;
wire _02896_;
wire _02897_;
wire _02898_;
wire _02899_;
wire _02900_;
wire _02901_;
wire _02902_;
wire _02903_;
wire _02904_;
wire _02905_;
wire _02906_;
wire _02907_;
wire _02908_;
wire _02909_;
wire _02910_;
wire _02911_;
wire _02912_;
wire _02913_;
wire _02914_;
wire _02915_;
wire _02916_;
wire _02917_;
wire _02918_;
wire _02919_;
wire _02920_;
wire _02921_;
wire _02922_;
wire _02923_;
wire _02924_;
wire _02925_;
wire _02926_;
wire _02927_;
wire _02928_;
wire _02929_;
wire _02930_;
wire _02931_;
wire _02932_;
wire _02933_;
wire _02934_;
wire _02935_;
wire _02936_;
wire _02937_;
wire _02938_;
wire _02939_;
wire _02940_;
wire _02941_;
wire _02942_;
wire _02943_;
wire _02944_;
wire _02945_;
wire _02946_;
wire _02947_;
wire _02948_;
wire _02949_;
wire _02950_;
wire _02951_;
wire _02952_;
wire _02953_;
wire _02954_;
wire _02955_;
wire _02956_;
wire _02957_;
wire _02958_;
wire _02959_;
wire _02960_;
wire _02961_;
wire _02962_;
wire _02963_;
wire _02964_;
wire _02965_;
wire _02966_;
wire _02967_;
wire _02968_;
wire _02969_;
wire _02970_;
wire _02971_;
wire _02972_;
wire _02973_;
wire _02974_;
wire _02975_;
wire _02976_;
wire _02977_;
wire _02978_;
wire _02979_;
wire _02980_;
wire _02981_;
wire _02982_;
wire _02983_;
wire _02984_;
wire _02985_;
wire _02986_;
wire _02987_;
wire _02988_;
wire _02989_;
wire _02990_;
wire _02991_;
wire _02992_;
wire _02993_;
wire _02994_;
wire _02995_;
wire _02996_;
wire _02997_;
wire _02998_;
wire _02999_;
wire _03000_;
wire _03001_;
wire _03002_;
wire _03003_;
wire _03004_;
wire _03005_;
wire _03006_;
wire _03007_;
wire _03008_;
wire _03009_;
wire _03010_;
wire _03011_;
wire _03012_;
wire _03013_;
wire _03014_;
wire _03015_;
wire _03016_;
wire _03017_;
wire _03018_;
wire _03019_;
wire _03020_;
wire _03021_;
wire _03022_;
wire _03023_;
wire _03024_;
wire _03025_;
wire _03026_;
wire _03027_;
wire _03028_;
wire _03029_;
wire _03030_;
wire _03031_;
wire _03032_;
wire _03033_;
wire _03034_;
wire _03035_;
wire _03036_;
wire _03037_;
wire _03038_;
wire _03039_;
wire _03040_;
wire _03041_;
wire _03042_;
wire _03043_;
wire _03044_;
wire _03045_;
wire _03046_;
wire _03047_;
wire _03048_;
wire _03049_;
wire _03050_;
wire _03051_;
wire _03052_;
wire _03053_;
wire _03054_;
wire _03055_;
wire _03056_;
wire _03057_;
wire _03058_;
wire _03059_;
wire _03060_;
wire _03061_;
wire _03062_;
wire _03063_;
wire _03064_;
wire _03065_;
wire _03066_;
wire _03067_;
wire _03068_;
wire _03069_;
wire _03070_;
wire _03071_;
wire _03072_;
wire _03073_;
wire _03074_;
wire _03075_;
wire _03076_;
wire _03077_;
wire _03078_;
wire _03079_;
wire _03080_;
wire _03081_;
wire _03082_;
wire _03083_;
wire _03084_;
wire _03085_;
wire _03086_;
wire _03087_;
wire _03088_;
wire _03089_;
wire _03090_;
wire _03091_;
wire _03092_;
wire _03093_;
wire _03094_;
wire _03095_;
wire _03096_;
wire _03097_;
wire _03098_;
wire _03099_;
wire _03100_;
wire _03101_;
wire _03102_;
wire _03103_;
wire _03104_;
wire _03105_;
wire _03106_;
wire _03107_;
wire _03108_;
wire _03109_;
wire _03110_;
wire _03111_;
wire _03112_;
wire _03113_;
wire _03114_;
wire _03115_;
wire _03116_;
wire _03117_;
wire _03118_;
wire _03119_;
wire _03120_;
wire _03121_;
wire _03122_;
wire _03123_;
wire _03124_;
wire _03125_;
wire _03126_;
wire _03127_;
wire _03128_;
wire _03129_;
wire _03130_;
wire _03131_;
wire _03132_;
wire _03133_;
wire _03134_;
wire _03135_;
wire _03136_;
wire _03137_;
wire _03138_;
wire _03139_;
wire _03140_;
wire _03141_;
wire _03142_;
wire _03143_;
wire _03144_;
wire _03145_;
wire _03146_;
wire _03147_;
wire _03148_;
wire _03149_;
wire _03150_;
wire _03151_;
wire _03152_;
wire _03153_;
wire _03154_;
wire _03155_;
wire _03156_;
wire _03157_;
wire _03158_;
wire _03159_;
wire _03160_;
wire _03161_;
wire _03162_;
wire _03163_;
wire _03164_;
wire _03165_;
wire _03166_;
wire _03167_;
wire _03168_;
wire _03169_;
wire _03170_;
wire _03171_;
wire _03172_;
wire _03173_;
wire _03174_;
wire _03175_;
wire _03176_;
wire _03177_;
wire _03178_;
wire _03179_;
wire _03180_;
wire _03181_;
wire _03182_;
wire _03183_;
wire _03184_;
wire _03185_;
wire _03186_;
wire _03187_;
wire _03188_;
wire _03189_;
wire _03190_;
wire _03191_;
wire _03192_;
wire _03193_;
wire _03194_;
wire _03195_;
wire _03196_;
wire _03197_;
wire _03198_;
wire _03199_;
wire _03200_;
wire _03201_;
wire _03202_;
wire _03203_;
wire _03204_;
wire _03205_;
wire _03206_;
wire _03207_;
wire _03208_;
wire _03209_;
wire _03210_;
wire _03211_;
wire _03212_;
wire _03213_;
wire _03214_;
wire _03215_;
wire _03216_;
wire _03217_;
wire _03218_;
wire _03219_;
wire _03220_;
wire _03221_;
wire _03222_;
wire _03223_;
wire _03224_;
wire _03225_;
wire _03226_;
wire _03227_;
wire _03228_;
wire _03229_;
wire _03230_;
wire _03231_;
wire _03232_;
wire _03233_;
wire _03234_;
wire _03235_;
wire _03236_;
wire _03237_;
wire _03238_;
wire _03239_;
wire _03240_;
wire _03241_;
wire _03242_;
wire _03243_;
wire _03244_;
wire _03245_;
wire _03246_;
wire _03247_;
wire _03248_;
wire _03249_;
wire _03250_;
wire _03251_;
wire _03252_;
wire _03253_;
wire _03254_;
wire _03255_;
wire _03256_;
wire _03257_;
wire _03258_;
wire _03259_;
wire _03260_;
wire _03261_;
wire _03262_;
wire _03263_;
wire _03264_;
wire _03265_;
wire _03266_;
wire _03267_;
wire _03268_;
wire _03269_;
wire _03270_;
wire _03271_;
wire _03272_;
wire _03273_;
wire _03274_;
wire _03275_;
wire _03276_;
wire _03277_;
wire _03278_;
wire _03279_;
wire _03280_;
wire _03281_;
wire _03282_;
wire _03283_;
wire _03284_;
wire _03285_;
wire _03286_;
wire _03287_;
wire _03288_;
wire _03289_;
wire _03290_;
wire _03291_;
wire _03292_;
wire _03293_;
wire _03294_;
wire _03295_;
wire _03296_;
wire _03297_;
wire _03298_;
wire _03299_;
wire _03300_;
wire _03301_;
wire _03302_;
wire _03303_;
wire _03304_;
wire _03305_;
wire _03306_;
wire _03307_;
wire _03308_;
wire _03309_;
wire _03310_;
wire _03311_;
wire _03312_;
wire _03313_;
wire _03314_;
wire _03315_;
wire _03316_;
wire _03317_;
wire _03318_;
wire _03319_;
wire _03320_;
wire _03321_;
wire _03322_;
wire _03323_;
wire _03324_;
wire _03325_;
wire _03326_;
wire _03327_;
wire _03328_;
wire _03329_;
wire _03330_;
wire _03331_;
wire _03332_;
wire _03333_;
wire _03334_;
wire _03335_;
wire _03336_;
wire _03337_;
wire _03338_;
wire _03339_;
wire _03340_;
wire _03341_;
wire _03342_;
wire _03343_;
wire _03344_;
wire _03345_;
wire _03346_;
wire _03347_;
wire _03348_;
wire _03349_;
wire _03350_;
wire _03351_;
wire _03352_;
wire _03353_;
wire _03354_;
wire _03355_;
wire _03356_;
wire _03357_;
wire _03358_;
wire _03359_;
wire _03360_;
wire _03361_;
wire _03362_;
wire _03363_;
wire _03364_;
wire _03365_;
wire _03366_;
wire _03367_;
wire _03368_;
wire _03369_;
wire _03370_;
wire _03371_;
wire _03372_;
wire _03373_;
wire _03374_;
wire _03375_;
wire _03376_;
wire _03377_;
wire _03378_;
wire _03379_;
wire _03380_;
wire _03381_;
wire _03382_;
wire _03383_;
wire _03384_;
wire _03385_;
wire _03386_;
wire _03387_;
wire _03388_;
wire _03389_;
wire _03390_;
wire _03391_;
wire _03392_;
wire _03393_;
wire _03394_;
wire _03395_;
wire _03396_;
wire _03397_;
wire _03398_;
wire _03399_;
wire _03400_;
wire _03401_;
wire _03402_;
wire _03403_;
wire _03404_;
wire _03405_;
wire _03406_;
wire _03407_;
wire _03408_;
wire _03409_;
wire _03410_;
wire _03411_;
wire _03412_;
wire _03413_;
wire _03414_;
wire _03415_;
wire _03416_;
wire _03417_;
wire _03418_;
wire _03419_;
wire _03420_;
wire _03421_;
wire _03422_;
wire _03423_;
wire _03424_;
wire _03425_;
wire _03426_;
wire _03427_;
wire _03428_;
wire _03429_;
wire _03430_;
wire _03431_;
wire _03432_;
wire _03433_;
wire _03434_;
wire _03435_;
wire _03436_;
wire _03437_;
wire _03438_;
wire _03439_;
wire _03440_;
wire _03441_;
wire _03442_;
wire _03443_;
wire _03444_;
wire _03445_;
wire _03446_;
wire _03447_;
wire _03448_;
wire _03449_;
wire _03450_;
wire _03451_;
wire _03452_;
wire _03453_;
wire _03454_;
wire _03455_;
wire _03456_;
wire _03457_;
wire _03458_;
wire _03459_;
wire _03460_;
wire _03461_;
wire _03462_;
wire _03463_;
wire _03464_;
wire _03465_;
wire _03466_;
wire _03467_;
wire _03468_;
wire _03469_;
wire _03470_;
wire _03471_;
wire _03472_;
wire _03473_;
wire _03474_;
wire _03475_;
wire _03476_;
wire _03477_;
wire _03478_;
wire _03479_;
wire _03480_;
wire _03481_;
wire _03482_;
wire _03483_;
wire _03484_;
wire _03485_;
wire _03486_;
wire _03487_;
wire _03488_;
wire _03489_;
wire _03490_;
wire _03491_;
wire _03492_;
wire _03493_;
wire _03494_;
wire _03495_;
wire _03496_;
wire _03497_;
wire _03498_;
wire _03499_;
wire _03500_;
wire _03501_;
wire _03502_;
wire _03503_;
wire _03504_;
wire _03505_;
wire _03506_;
wire _03507_;
wire _03508_;
wire _03509_;
wire _03510_;
wire _03511_;
wire _03512_;
wire _03513_;
wire _03514_;
wire _03515_;
wire _03516_;
wire _03517_;
wire _03518_;
wire _03519_;
wire _03520_;
wire _03521_;
wire _03522_;
wire _03523_;
wire _03524_;
wire _03525_;
wire _03526_;
wire _03527_;
wire _03528_;
wire _03529_;
wire _03530_;
wire _03531_;
wire _03532_;
wire _03533_;
wire _03534_;
wire _03535_;
wire _03536_;
wire _03537_;
wire _03538_;
wire _03539_;
wire _03540_;
wire _03541_;
wire _03542_;
wire _03543_;
wire _03544_;
wire _03545_;
wire _03546_;
wire _03547_;
wire _03548_;
wire _03549_;
wire _03550_;
wire _03551_;
wire _03552_;
wire _03553_;
wire _03554_;
wire _03555_;
wire _03556_;
wire _03557_;
wire _03558_;
wire _03559_;
wire _03560_;
wire _03561_;
wire _03562_;
wire _03563_;
wire _03564_;
wire _03565_;
wire _03566_;
wire _03567_;
wire _03568_;
wire _03569_;
wire _03570_;
wire _03571_;
wire _03572_;
wire _03573_;
wire _03574_;
wire _03575_;
wire _03576_;
wire _03577_;
wire _03578_;
wire _03579_;
wire _03580_;
wire _03581_;
wire _03582_;
wire _03583_;
wire _03584_;
wire _03585_;
wire _03586_;
wire _03587_;
wire _03588_;
wire _03589_;
wire _03590_;
wire _03591_;
wire _03592_;
wire _03593_;
wire _03594_;
wire _03595_;
wire _03596_;
wire _03597_;
wire _03598_;
wire _03599_;
wire _03600_;
wire _03601_;
wire _03602_;
wire _03603_;
wire _03604_;
wire _03605_;
wire _03606_;
wire _03607_;
wire _03608_;
wire _03609_;
wire _03610_;
wire _03611_;
wire _03612_;
wire _03613_;
wire _03614_;
wire _03615_;
wire _03616_;
wire _03617_;
wire _03618_;
wire _03619_;
wire _03620_;
wire _03621_;
wire _03622_;
wire _03623_;
wire _03624_;
wire _03625_;
wire _03626_;
wire _03627_;
wire _03628_;
wire _03629_;
wire _03630_;
wire _03631_;
wire _03632_;
wire _03633_;
wire _03634_;
wire _03635_;
wire _03636_;
wire _03637_;
wire _03638_;
wire _03639_;
wire _03640_;
wire _03641_;
wire _03642_;
wire _03643_;
wire _03644_;
wire _03645_;
wire _03646_;
wire _03647_;
wire _03648_;
wire _03649_;
wire _03650_;
wire _03651_;
wire _03652_;
wire _03653_;
wire _03654_;
wire _03655_;
wire _03656_;
wire _03657_;
wire _03658_;
wire _03659_;
wire _03660_;
wire _03661_;
wire _03662_;
wire _03663_;
wire _03664_;
wire _03665_;
wire _03666_;
wire _03667_;
wire _03668_;
wire _03669_;
wire _03670_;
wire _03671_;
wire _03672_;
wire _03673_;
wire _03674_;
wire _03675_;
wire _03676_;
wire _03677_;
wire _03678_;
wire _03679_;
wire _03680_;
wire _03681_;
wire _03682_;
wire _03683_;
wire _03684_;
wire _03685_;
wire _03686_;
wire _03687_;
wire _03688_;
wire _03689_;
wire _03690_;
wire _03691_;
wire _03692_;
wire _03693_;
wire _03694_;
wire _03695_;
wire _03696_;
wire _03697_;
wire _03698_;
wire _03699_;
wire _03700_;
wire _03701_;
wire _03702_;
wire _03703_;
wire _03704_;
wire _03705_;
wire _03706_;
wire _03707_;
wire _03708_;
wire _03709_;
wire _03710_;
wire _03711_;
wire _03712_;
wire _03713_;
wire _03714_;
wire _03715_;
wire _03716_;
wire _03717_;
wire _03718_;
wire _03719_;
wire _03720_;
wire _03721_;
wire _03722_;
wire _03723_;
wire _03724_;
wire _03725_;
wire _03726_;
wire _03727_;
wire _03728_;
wire _03729_;
wire _03730_;
wire _03731_;
wire _03732_;
wire _03733_;
wire _03734_;
wire _03735_;
wire _03736_;
wire _03737_;
wire _03738_;
wire _03739_;
wire _03740_;
wire _03741_;
wire _03742_;
wire _03743_;
wire _03744_;
wire _03745_;
wire _03746_;
wire _03747_;
wire _03748_;
wire _03749_;
wire _03750_;
wire _03751_;
wire _03752_;
wire _03753_;
wire _03754_;
wire _03755_;
wire _03756_;
wire _03757_;
wire _03758_;
wire _03759_;
wire _03760_;
wire _03761_;
wire _03762_;
wire _03763_;
wire _03764_;
wire _03765_;
wire _03766_;
wire _03767_;
wire _03768_;
wire _03769_;
wire _03770_;
wire _03771_;
wire _03772_;
wire _03773_;
wire _03774_;
wire _03775_;
wire _03776_;
wire _03777_;
wire _03778_;
wire _03779_;
wire _03780_;
wire _03781_;
wire _03782_;
wire _03783_;
wire _03784_;
wire _03785_;
wire _03786_;
wire _03787_;
wire _03788_;
wire _03789_;
wire _03790_;
wire _03791_;
wire _03792_;
wire _03793_;
wire _03794_;
wire _03795_;
wire _03796_;
wire _03797_;
wire _03798_;
wire _03799_;
wire _03800_;
wire _03801_;
wire _03802_;
wire _03803_;
wire _03804_;
wire _03805_;
wire _03806_;
wire _03807_;
wire _03808_;
wire _03809_;
wire _03810_;
wire _03811_;
wire _03812_;
wire _03813_;
wire _03814_;
wire _03815_;
wire _03816_;
wire _03817_;
wire _03818_;
wire _03819_;
wire _03820_;
wire _03821_;
wire _03822_;
wire _03823_;
wire _03824_;
wire _03825_;
wire _03826_;
wire _03827_;
wire _03828_;
wire _03829_;
wire _03830_;
wire _03831_;
wire _03832_;
wire _03833_;
wire _03834_;
wire _03835_;
wire _03836_;
wire _03837_;
wire _03838_;
wire _03839_;
wire _03840_;
wire _03841_;
wire _03842_;
wire _03843_;
wire _03844_;
wire _03845_;
wire _03846_;
wire _03847_;
wire _03848_;
wire _03849_;
wire _03850_;
wire _03851_;
wire _03852_;
wire _03853_;
wire _03854_;
wire _03855_;
wire _03856_;
wire _03857_;
wire _03858_;
wire _03859_;
wire _03860_;
wire _03861_;
wire _03862_;
wire _03863_;
wire _03864_;
wire _03865_;
wire _03866_;
wire _03867_;
wire _03868_;
wire _03869_;
wire _03870_;
wire _03871_;
wire _03872_;
wire _03873_;
wire _03874_;
wire _03875_;
wire _03876_;
wire _03877_;
wire _03878_;
wire _03879_;
wire _03880_;
wire _03881_;
wire _03882_;
wire _03883_;
wire _03884_;
wire _03885_;
wire _03886_;
wire _03887_;
wire _03888_;
wire _03889_;
wire _03890_;
wire _03891_;
wire _03892_;
wire _03893_;
wire _03894_;
wire _03895_;
wire _03896_;
wire _03897_;
wire _03898_;
wire _03899_;
wire _03900_;
wire _03901_;
wire _03902_;
wire _03903_;
wire _03904_;
wire _03905_;
wire _03906_;
wire _03907_;
wire _03908_;
wire _03909_;
wire _03910_;
wire _03911_;
wire _03912_;
wire _03913_;
wire _03914_;
wire _03915_;
wire _03916_;
wire _03917_;
wire _03918_;
wire _03919_;
wire _03920_;
wire _03921_;
wire _03922_;
wire _03923_;
wire _03924_;
wire _03925_;
wire _03926_;
wire _03927_;
wire _03928_;
wire _03929_;
wire _03930_;
wire _03931_;
wire _03932_;
wire _03933_;
wire _03934_;
wire _03935_;
wire _03936_;
wire _03937_;
wire _03938_;
wire _03939_;
wire _03940_;
wire _03941_;
wire _03942_;
wire _03943_;
wire _03944_;
wire _03945_;
wire _03946_;
wire _03947_;
wire _03948_;
wire _03949_;
wire _03950_;
wire _03951_;
wire _03952_;
wire _03953_;
wire _03954_;
wire _03955_;
wire _03956_;
wire _03957_;
wire _03958_;
wire _03959_;
wire _03960_;
wire _03961_;
wire _03962_;
wire _03963_;
wire _03964_;
wire _03965_;
wire _03966_;
wire _03967_;
wire _03968_;
wire _03969_;
wire _03970_;
wire _03971_;
wire _03972_;
wire _03973_;
wire _03974_;
wire _03975_;
wire _03976_;
wire _03977_;
wire _03978_;
wire _03979_;
wire _03980_;
wire _03981_;
wire _03982_;
wire _03983_;
wire _03984_;
wire _03985_;
wire _03986_;
wire _03987_;
wire _03988_;
wire _03989_;
wire _03990_;
wire _03991_;
wire _03992_;
wire _03993_;
wire _03994_;
wire _03995_;
wire _03996_;
wire _03997_;
wire _03998_;
wire _03999_;
wire _04000_;
wire _04001_;
wire _04002_;
wire _04003_;
wire _04004_;
wire _04005_;
wire _04006_;
wire _04007_;
wire _04008_;
wire _04009_;
wire _04010_;
wire _04011_;
wire _04012_;
wire _04013_;
wire _04014_;
wire _04015_;
wire _04016_;
wire _04017_;
wire _04018_;
wire _04019_;
wire _04020_;
wire _04021_;
wire _04022_;
wire _04023_;
wire _04024_;
wire _04025_;
wire _04026_;
wire _04027_;
wire _04028_;
wire _04029_;
wire _04030_;
wire _04031_;
wire _04032_;
wire _04033_;
wire _04034_;
wire _04035_;
wire _04036_;
wire _04037_;
wire _04038_;
wire _04039_;
wire _04040_;
wire _04041_;
wire _04042_;
wire _04043_;
wire _04044_;
wire _04045_;
wire _04046_;
wire _04047_;
wire _04048_;
wire _04049_;
wire _04050_;
wire _04051_;
wire _04052_;
wire _04053_;
wire _04054_;
wire _04055_;
wire _04056_;
wire _04057_;
wire _04058_;
wire _04059_;
wire _04060_;
wire _04061_;
wire _04062_;
wire _04063_;
wire _04064_;
wire _04065_;
wire _04066_;
wire _04067_;
wire _04068_;
wire _04069_;
wire _04070_;
wire _04071_;
wire _04072_;
wire _04073_;
wire _04074_;
wire _04075_;
wire _04076_;
wire _04077_;
wire _04078_;
wire _04079_;
wire _04080_;
wire _04081_;
wire _04082_;
wire _04083_;
wire _04084_;
wire _04085_;
wire _04086_;
wire _04087_;
wire _04088_;
wire _04089_;
wire _04090_;
wire _04091_;
wire _04092_;
wire _04093_;
wire _04094_;
wire _04095_;
wire _04096_;
wire _04097_;
wire _04098_;
wire _04099_;
wire _04100_;
wire _04101_;
wire _04102_;
wire _04103_;
wire _04104_;
wire _04105_;
wire _04106_;
wire _04107_;
wire _04108_;
wire _04109_;
wire _04110_;
wire _04111_;
wire _04112_;
wire _04113_;
wire _04114_;
wire _04115_;
wire _04116_;
wire _04117_;
wire _04118_;
wire _04119_;
wire _04120_;
wire _04121_;
wire _04122_;
wire _04123_;
wire _04124_;
wire _04125_;
wire _04126_;
wire _04127_;
wire _04128_;
wire _04129_;
wire _04130_;
wire _04131_;
wire _04132_;
wire _04133_;
wire _04134_;
wire _04135_;
wire _04136_;
wire _04137_;
wire _04138_;
wire _04139_;
wire _04140_;
wire _04141_;
wire _04142_;
wire _04143_;
wire _04144_;
wire _04145_;
wire _04146_;
wire _04147_;
wire _04148_;
wire _04149_;
wire _04150_;
wire _04151_;
wire _04152_;
wire _04153_;
wire _04154_;
wire _04155_;
wire _04156_;
wire _04157_;
wire _04158_;
wire _04159_;
wire _04160_;
wire _04161_;
wire _04162_;
wire _04163_;
wire _04164_;
wire _04165_;
wire _04166_;
wire _04167_;
wire _04168_;
wire _04169_;
wire _04170_;
wire _04171_;
wire _04172_;
wire _04173_;
wire _04174_;
wire _04175_;
wire _04176_;
wire _04177_;
wire _04178_;
wire _04179_;
wire _04180_;
wire _04181_;
wire _04182_;
wire _04183_;
wire _04184_;
wire _04185_;
wire _04186_;
wire _04187_;
wire _04188_;
wire _04189_;
wire _04190_;
wire _04191_;
wire _04192_;
wire _04193_;
wire _04194_;
wire _04195_;
wire _04196_;
wire _04197_;
wire _04198_;
wire _04199_;
wire _04200_;
wire _04201_;
wire _04202_;
wire _04203_;
wire _04204_;
wire _04205_;
wire _04206_;
wire _04207_;
wire _04208_;
wire _04209_;
wire _04210_;
wire _04211_;
wire _04212_;
wire _04213_;
wire _04214_;
wire _04215_;
wire _04216_;
wire _04217_;
wire _04218_;
wire _04219_;
wire _04220_;
wire _04221_;
wire _04222_;
wire _04223_;
wire _04224_;
wire _04225_;
wire _04226_;
wire _04227_;
wire _04228_;
wire _04229_;
wire _04230_;
wire _04231_;
wire _04232_;
wire _04233_;
wire _04234_;
wire _04235_;
wire _04236_;
wire _04237_;
wire _04238_;
wire _04239_;
wire _04240_;
wire _04241_;
wire _04242_;
wire _04243_;
wire _04244_;
wire _04245_;
wire _04246_;
wire _04247_;
wire _04248_;
wire _04249_;
wire _04250_;
wire _04251_;
wire _04252_;
wire _04253_;
wire _04254_;
wire _04255_;
wire _04256_;
wire _04257_;
wire _04258_;
wire _04259_;
wire _04260_;
wire _04261_;
wire _04262_;
wire _04263_;
wire _04264_;
wire _04265_;
wire _04266_;
wire _04267_;
wire _04268_;
wire _04269_;
wire _04270_;
wire _04271_;
wire _04272_;
wire _04273_;
wire _04274_;
wire _04275_;
wire _04276_;
wire _04277_;
wire _04278_;
wire _04279_;
wire _04280_;
wire _04281_;
wire _04282_;
wire _04283_;
wire _04284_;
wire _04285_;
wire _04286_;
wire _04287_;
wire _04288_;
wire _04289_;
wire _04290_;
wire _04291_;
wire _04292_;
wire _04293_;
wire _04294_;
wire _04295_;
wire _04296_;
wire _04297_;
wire _04298_;
wire _04299_;
wire _04300_;
wire _04301_;
wire _04302_;
wire _04303_;
wire _04304_;
wire _04305_;
wire _04306_;
wire _04307_;
wire _04308_;
wire _04309_;
wire _04310_;
wire _04311_;
wire _04312_;
wire _04313_;
wire _04314_;
wire _04315_;
wire _04316_;
wire _04317_;
wire _04318_;
wire _04319_;
wire _04320_;
wire _04321_;
wire _04322_;
wire _04323_;
wire _04324_;
wire _04325_;
wire _04326_;
wire _04327_;
wire _04328_;
wire _04329_;
wire _04330_;
wire _04331_;
wire _04332_;
wire _04333_;
wire _04334_;
wire _04335_;
wire _04336_;
wire _04337_;
wire _04338_;
wire _04339_;
wire _04340_;
wire _04341_;
wire _04342_;
wire _04343_;
wire _04344_;
wire _04345_;
wire _04346_;
wire _04347_;
wire _04348_;
wire _04349_;
wire _04350_;
wire _04351_;
wire _04352_;
wire _04353_;
wire _04354_;
wire _04355_;
wire _04356_;
wire _04357_;
wire _04358_;
wire _04359_;
wire _04360_;
wire _04361_;
wire _04362_;
wire _04363_;
wire _04364_;
wire _04365_;
wire _04366_;
wire _04367_;
wire _04368_;
wire _04369_;
wire _04370_;
wire _04371_;
wire _04372_;
wire _04373_;
wire _04374_;
wire _04375_;
wire _04376_;
wire _04377_;
wire _04378_;
wire _04379_;
wire _04380_;
wire _04381_;
wire _04382_;
wire _04383_;
wire _04384_;
wire _04385_;
wire _04386_;
wire _04387_;
wire _04388_;
wire _04389_;
wire _04390_;
wire _04391_;
wire _04392_;
wire _04393_;
wire _04394_;
wire _04395_;
wire _04396_;
wire _04397_;
wire _04398_;
wire _04399_;
wire _04400_;
wire _04401_;
wire _04402_;
wire _04403_;
wire _04404_;
wire _04405_;
wire _04406_;
wire _04407_;
wire _04408_;
wire _04409_;
wire _04410_;
wire _04411_;
wire _04412_;
wire _04413_;
wire _04414_;
wire _04415_;
wire _04416_;
wire _04417_;
wire _04418_;
wire _04419_;
wire _04420_;
wire _04421_;
wire _04422_;
wire _04423_;
wire _04424_;
wire _04425_;
wire _04426_;
wire _04427_;
wire _04428_;
wire _04429_;
wire _04430_;
wire _04431_;
wire _04432_;
wire _04433_;
wire _04434_;
wire _04435_;
wire _04436_;
wire _04437_;
wire _04438_;
wire _04439_;
wire _04440_;
wire _04441_;
wire _04442_;
wire _04443_;
wire _04444_;
wire _04445_;
wire _04446_;
wire _04447_;
wire _04448_;
wire _04449_;
wire _04450_;
wire _04451_;
wire _04452_;
wire _04453_;
wire _04454_;
wire _04455_;
wire _04456_;
wire _04457_;
wire _04458_;
wire _04459_;
wire _04460_;
wire _04461_;
wire _04462_;
wire _04463_;
wire _04464_;
wire _04465_;
wire _04466_;
wire _04467_;
wire _04468_;
wire _04469_;
wire _04470_;
wire _04471_;
wire _04472_;
wire _04473_;
wire _04474_;
wire _04475_;
wire _04476_;
wire _04477_;
wire _04478_;
wire _04479_;
wire _04480_;
wire _04481_;
wire _04482_;
wire _04483_;
wire _04484_;
wire _04485_;
wire _04486_;
wire _04487_;
wire _04488_;
wire _04489_;
wire _04490_;
wire _04491_;
wire _04492_;
wire _04493_;
wire _04494_;
wire _04495_;
wire _04496_;
wire _04497_;
wire _04498_;
wire _04499_;
wire _04500_;
wire _04501_;
wire _04502_;
wire _04503_;
wire _04504_;
wire _04505_;
wire _04506_;
wire _04507_;
wire _04508_;
wire _04509_;
wire _04510_;
wire _04511_;
wire _04512_;
wire _04513_;
wire _04514_;
wire _04515_;
wire _04516_;
wire _04517_;
wire _04518_;
wire _04519_;
wire _04520_;
wire _04521_;
wire _04522_;
wire _04523_;
wire _04524_;
wire _04525_;
wire _04526_;
wire _04527_;
wire _04528_;
wire _04529_;
wire _04530_;
wire _04531_;
wire _04532_;
wire _04533_;
wire _04534_;
wire _04535_;
wire _04536_;
wire _04537_;
wire _04538_;
wire _04539_;
wire _04540_;
wire _04541_;
wire _04542_;
wire _04543_;
wire _04544_;
wire _04545_;
wire _04546_;
wire _04547_;
wire _04548_;
wire _04549_;
wire _04550_;
wire _04551_;
wire _04552_;
wire _04553_;
wire _04554_;
wire _04555_;
wire _04556_;
wire _04557_;
wire _04558_;
wire _04559_;
wire _04560_;
wire _04561_;
wire _04562_;
wire _04563_;
wire _04564_;
wire _04565_;
wire _04566_;
wire _04567_;
wire _04568_;
wire _04569_;
wire _04570_;
wire _04571_;
wire _04572_;
wire _04573_;
wire _04574_;
wire _04575_;
wire _04576_;
wire _04577_;
wire _04578_;
wire _04579_;
wire _04580_;
wire _04581_;
wire _04582_;
wire _04583_;
wire _04584_;
wire _04585_;
wire _04586_;
wire _04587_;
wire _04588_;
wire _04589_;
wire _04590_;
wire _04591_;
wire _04592_;
wire _04593_;
wire _04594_;
wire _04595_;
wire _04596_;
wire _04597_;
wire _04598_;
wire _04599_;
wire _04600_;
wire _04601_;
wire _04602_;
wire _04603_;
wire _04604_;
wire _04605_;
wire _04606_;
wire _04607_;
wire _04608_;
wire _04609_;
wire _04610_;
wire _04611_;
wire _04612_;
wire _04613_;
wire _04614_;
wire _04615_;
wire _04616_;
wire _04617_;
wire _04618_;
wire _04619_;
wire _04620_;
wire _04621_;
wire _04622_;
wire _04623_;
wire _04624_;
wire _04625_;
wire _04626_;
wire _04627_;
wire _04628_;
wire _04629_;
wire _04630_;
wire _04631_;
wire _04632_;
wire _04633_;
wire _04634_;
wire _04635_;
wire _04636_;
wire _04637_;
wire _04638_;
wire _04639_;
wire _04640_;
wire _04641_;
wire _04642_;
wire _04643_;
wire _04644_;
wire _04645_;
wire _04646_;
wire _04647_;
wire _04648_;
wire _04649_;
wire _04650_;
wire _04651_;
wire _04652_;
wire _04653_;
wire _04654_;
wire _04655_;
wire _04656_;
wire _04657_;
wire _04658_;
wire _04659_;
wire _04660_;
wire _04661_;
wire _04662_;
wire _04663_;
wire _04664_;
wire _04665_;
wire _04666_;
wire _04667_;
wire _04668_;
wire _04669_;
wire _04670_;
wire _04671_;
wire _04672_;
wire _04673_;
wire _04674_;
wire _04675_;
wire _04676_;
wire _04677_;
wire _04678_;
wire _04679_;
wire _04680_;
wire _04681_;
wire _04682_;
wire _04683_;
wire _04684_;
wire _04685_;
wire _04686_;
wire _04687_;
wire _04688_;
wire _04689_;
wire _04690_;
wire _04691_;
wire _04692_;
wire _04693_;
wire _04694_;
wire _04695_;
wire _04696_;
wire _04697_;
wire _04698_;
wire _04699_;
wire _04700_;
wire _04701_;
wire _04702_;
wire _04703_;
wire _04704_;
wire _04705_;
wire _04706_;
wire _04707_;
wire _04708_;
wire _04709_;
wire _04710_;
wire _04711_;
wire _04712_;
wire _04713_;
wire _04714_;
wire _04715_;
wire _04716_;
wire _04717_;
wire _04718_;
wire _04719_;
wire _04720_;
wire _04721_;
wire _04722_;
wire _04723_;
wire _04724_;
wire _04725_;
wire _04726_;
wire _04727_;
wire _04728_;
wire _04729_;
wire _04730_;
wire _04731_;
wire _04732_;
wire _04733_;
wire _04734_;
wire _04735_;
wire _04736_;
wire _04737_;
wire _04738_;
wire _04739_;
wire _04740_;
wire _04741_;
wire _04742_;
wire _04743_;
wire _04744_;
wire _04745_;
wire _04746_;
wire _04747_;
wire _04748_;
wire _04749_;
wire _04750_;
wire _04751_;
wire _04752_;
wire _04753_;
wire _04754_;
wire _04755_;
wire _04756_;
wire _04757_;
wire _04758_;
wire _04759_;
wire _04760_;
wire _04761_;
wire _04762_;
wire _04763_;
wire _04764_;
wire _04765_;
wire _04766_;
wire _04767_;
wire _04768_;
wire _04769_;
wire _04770_;
wire _04771_;
wire _04772_;
wire _04773_;
wire _04774_;
wire _04775_;
wire _04776_;
wire _04777_;
wire _04778_;
wire _04779_;
wire _04780_;
wire _04781_;
wire _04782_;
wire _04783_;
wire _04784_;
wire _04785_;
wire _04786_;
wire _04787_;
wire _04788_;
wire _04789_;
wire _04790_;
wire _04791_;
wire _04792_;
wire _04793_;
wire _04794_;
wire _04795_;
wire _04796_;
wire _04797_;
wire _04798_;
wire _04799_;
wire _04800_;
wire _04801_;
wire _04802_;
wire _04803_;
wire _04804_;
wire _04805_;
wire _04806_;
wire _04807_;
wire _04808_;
wire _04809_;
wire _04810_;
wire _04811_;
wire _04812_;
wire _04813_;
wire _04814_;
wire _04815_;
wire _04816_;
wire _04817_;
wire _04818_;
wire _04819_;
wire _04820_;
wire _04821_;
wire _04822_;
wire _04823_;
wire _04824_;
wire _04825_;
wire _04826_;
wire _04827_;
wire _04828_;
wire _04829_;
wire _04830_;
wire _04831_;
wire _04832_;
wire _04833_;
wire _04834_;
wire _04835_;
wire _04836_;
wire _04837_;
wire _04838_;
wire _04839_;
wire _04840_;
wire _04841_;
wire _04842_;
wire _04843_;
wire _04844_;
wire _04845_;
wire _04846_;
wire _04847_;
wire _04848_;
wire _04849_;
wire _04850_;
wire _04851_;
wire _04852_;
wire _04853_;
wire _04854_;
wire _04855_;
wire _04856_;
wire _04857_;
wire _04858_;
wire _04859_;
wire _04860_;
wire _04861_;
wire _04862_;
wire _04863_;
wire _04864_;
wire _04865_;
wire _04866_;
wire _04867_;
wire _04868_;
wire _04869_;
wire _04870_;
wire _04871_;
wire _04872_;
wire _04873_;
wire _04874_;
wire _04875_;
wire _04876_;
wire _04877_;
wire _04878_;
wire _04879_;
wire _04880_;
wire _04881_;
wire _04882_;
wire _04883_;
wire _04884_;
wire _04885_;
wire _04886_;
wire _04887_;
wire _04888_;
wire _04889_;
wire _04890_;
wire _04891_;
wire _04892_;
wire _04893_;
wire _04894_;
wire _04895_;
wire _04896_;
wire _04897_;
wire _04898_;
wire _04899_;
wire _04900_;
wire _04901_;
wire _04902_;
wire _04903_;
wire _04904_;
wire _04905_;
wire _04906_;
wire _04907_;
wire _04908_;
wire _04909_;
wire _04910_;
wire _04911_;
wire _04912_;
wire _04913_;
wire _04914_;
wire _04915_;
wire _04916_;
wire _04917_;
wire _04918_;
wire _04919_;
wire _04920_;
wire _04921_;
wire _04922_;
wire _04923_;
wire _04924_;
wire _04925_;
wire _04926_;
wire _04927_;
wire _04928_;
wire _04929_;
wire _04930_;
wire _04931_;
wire _04932_;
wire _04933_;
wire _04934_;
wire _04935_;
wire _04936_;
wire _04937_;
wire _04938_;
wire _04939_;
wire _04940_;
wire _04941_;
wire _04942_;
wire _04943_;
wire _04944_;
wire _04945_;
wire _04946_;
wire _04947_;
wire _04948_;
wire _04949_;
wire _04950_;
wire _04951_;
wire _04952_;
wire _04953_;
wire _04954_;
wire _04955_;
wire _04956_;
wire _04957_;
wire _04958_;
wire _04959_;
wire _04960_;
wire _04961_;
wire _04962_;
wire _04963_;
wire _04964_;
wire _04965_;
wire _04966_;
wire _04967_;
wire _04968_;
wire _04969_;
wire _04970_;
wire _04971_;
wire _04972_;
wire _04973_;
wire _04974_;
wire _04975_;
wire _04976_;
wire _04977_;
wire _04978_;
wire _04979_;
wire _04980_;
wire _04981_;
wire _04982_;
wire _04983_;
wire _04984_;
wire _04985_;
wire _04986_;
wire _04987_;
wire _04988_;
wire _04989_;
wire _04990_;
wire _04991_;
wire _04992_;
wire _04993_;
wire _04994_;
wire _04995_;
wire _04996_;
wire _04997_;
wire _04998_;
wire _04999_;
wire _05000_;
wire _05001_;
wire _05002_;
wire _05003_;
wire _05004_;
wire _05005_;
wire _05006_;
wire _05007_;
wire _05008_;
wire _05009_;
wire _05010_;
wire _05011_;
wire _05012_;
wire _05013_;
wire _05014_;
wire _05015_;
wire _05016_;
wire _05017_;
wire _05018_;
wire _05019_;
wire _05020_;
wire _05021_;
wire _05022_;
wire _05023_;
wire _05024_;
wire _05025_;
wire _05026_;
wire _05027_;
wire _05028_;
wire _05029_;
wire _05030_;
wire _05031_;
wire _05032_;
wire _05033_;
wire _05034_;
wire _05035_;
wire _05036_;
wire _05037_;
wire _05038_;
wire _05039_;
wire _05040_;
wire _05041_;
wire _05042_;
wire _05043_;
wire _05044_;
wire _05045_;
wire _05046_;
wire _05047_;
wire _05048_;
wire _05049_;
wire _05050_;
wire _05051_;
wire _05052_;
wire _05053_;
wire _05054_;
wire _05055_;
wire _05056_;
wire _05057_;
wire _05058_;
wire _05059_;
wire _05060_;
wire _05061_;
wire _05062_;
wire _05063_;
wire _05064_;
wire _05065_;
wire _05066_;
wire _05067_;
wire _05068_;
wire _05069_;
wire _05070_;
wire _05071_;
wire _05072_;
wire _05073_;
wire _05074_;
wire _05075_;
wire _05076_;
wire _05077_;
wire _05078_;
wire _05079_;
wire _05080_;
wire _05081_;
wire _05082_;
wire _05083_;
wire _05084_;
wire _05085_;
wire _05086_;
wire _05087_;
wire _05088_;
wire _05089_;
wire _05090_;
wire _05091_;
wire _05092_;
wire _05093_;
wire _05094_;
wire _05095_;
wire _05096_;
wire _05097_;
wire _05098_;
wire _05099_;
wire _05100_;
wire _05101_;
wire _05102_;
wire _05103_;
wire _05104_;
wire _05105_;
wire _05106_;
wire _05107_;
wire _05108_;
wire _05109_;
wire _05110_;
wire _05111_;
wire _05112_;
wire _05113_;
wire _05114_;
wire _05115_;
wire _05116_;
wire _05117_;
wire _05118_;
wire _05119_;
wire _05120_;
wire _05121_;
wire _05122_;
wire _05123_;
wire _05124_;
wire _05125_;
wire _05126_;
wire _05127_;
wire _05128_;
wire _05129_;
wire _05130_;
wire _05131_;
wire _05132_;
wire _05133_;
wire _05134_;
wire _05135_;
wire _05136_;
wire _05137_;
wire _05138_;
wire _05139_;
wire _05140_;
wire _05141_;
wire _05142_;
wire _05143_;
wire _05144_;
wire _05145_;
wire _05146_;
wire _05147_;
wire _05148_;
wire _05149_;
wire _05150_;
wire _05151_;
wire _05152_;
wire _05153_;
wire _05154_;
wire _05155_;
wire _05156_;
wire _05157_;
wire _05158_;
wire _05159_;
wire _05160_;
wire _05161_;
wire _05162_;
wire _05163_;
wire _05164_;
wire _05165_;
wire _05166_;
wire _05167_;
wire _05168_;
wire _05169_;
wire _05170_;
wire _05171_;
wire _05172_;
wire _05173_;
wire _05174_;
wire _05175_;
wire _05176_;
wire _05177_;
wire _05178_;
wire _05179_;
wire _05180_;
wire _05181_;
wire _05182_;
wire _05183_;
wire _05184_;
wire _05185_;
wire _05186_;
wire _05187_;
wire _05188_;
wire _05189_;
wire _05190_;
wire _05191_;
wire _05192_;
wire _05193_;
wire _05194_;
wire _05195_;
wire _05196_;
wire _05197_;
wire _05198_;
wire _05199_;
wire _05200_;
wire _05201_;
wire _05202_;
wire _05203_;
wire _05204_;
wire _05205_;
wire _05206_;
wire _05207_;
wire _05208_;
wire _05209_;
wire _05210_;
wire _05211_;
wire _05212_;
wire _05213_;
wire _05214_;
wire _05215_;
wire _05216_;
wire _05217_;
wire _05218_;
wire _05219_;
wire _05220_;
wire _05221_;
wire _05222_;
wire _05223_;
wire _05224_;
wire _05225_;
wire _05226_;
wire _05227_;
wire _05228_;
wire _05229_;
wire _05230_;
wire _05231_;
wire _05232_;
wire _05233_;
wire _05234_;
wire _05235_;
wire _05236_;
wire _05237_;
wire _05238_;
wire _05239_;
wire _05240_;
wire _05241_;
wire _05242_;
wire _05243_;
wire _05244_;
wire _05245_;
wire _05246_;
wire _05247_;
wire _05248_;
wire _05249_;
wire _05250_;
wire _05251_;
wire _05252_;
wire _05253_;
wire _05254_;
wire _05255_;
wire _05256_;
wire _05257_;
wire _05258_;
wire _05259_;
wire _05260_;
wire _05261_;
wire _05262_;
wire _05263_;
wire _05264_;
wire _05265_;
wire _05266_;
wire _05267_;
wire _05268_;
wire _05269_;
wire _05270_;
wire _05271_;
wire _05272_;
wire _05273_;
wire _05274_;
wire _05275_;
wire _05276_;
wire _05277_;
wire _05278_;
wire _05279_;
wire _05280_;
wire _05281_;
wire _05282_;
wire _05283_;
wire _05284_;
wire _05285_;
wire _05286_;
wire _05287_;
wire _05288_;
wire _05289_;
wire _05290_;
wire _05291_;
wire _05292_;
wire _05293_;
wire _05294_;
wire _05295_;
wire _05296_;
wire _05297_;
wire _05298_;
wire _05299_;
wire _05300_;
wire _05301_;
wire _05302_;
wire _05303_;
wire _05304_;
wire _05305_;
wire _05306_;
wire _05307_;
wire _05308_;
wire _05309_;
wire _05310_;
wire _05311_;
wire _05312_;
wire _05313_;
wire _05314_;
wire _05315_;
wire _05316_;
wire _05317_;
wire _05318_;
wire _05319_;
wire _05320_;
wire _05321_;
wire _05322_;
wire _05323_;
wire _05324_;
wire _05325_;
wire _05326_;
wire _05327_;
wire _05328_;
wire _05329_;
wire _05330_;
wire _05331_;
wire _05332_;
wire _05333_;
wire _05334_;
wire _05335_;
wire _05336_;
wire _05337_;
wire _05338_;
wire _05339_;
wire _05340_;
wire _05341_;
wire _05342_;
wire _05343_;
wire _05344_;
wire _05345_;
wire _05346_;
wire _05347_;
wire _05348_;
wire _05349_;
wire _05350_;
wire _05351_;
wire _05352_;
wire _05353_;
wire _05354_;
wire _05355_;
wire _05356_;
wire _05357_;
wire _05358_;
wire _05359_;
wire _05360_;
wire _05361_;
wire _05362_;
wire _05363_;
wire _05364_;
wire _05365_;
wire _05366_;
wire _05367_;
wire _05368_;
wire _05369_;
wire _05370_;
wire _05371_;
wire _05372_;
wire _05373_;
wire _05374_;
wire _05375_;
wire _05376_;
wire _05377_;
wire _05378_;
wire _05379_;
wire _05380_;
wire _05381_;
wire _05382_;
wire _05383_;
wire _05384_;
wire _05385_;
wire _05386_;
wire _05387_;
wire _05388_;
wire _05389_;
wire _05390_;
wire _05391_;
wire _05392_;
wire _05393_;
wire _05394_;
wire _05395_;
wire _05396_;
wire _05397_;
wire _05398_;
wire _05399_;
wire _05400_;
wire _05401_;
wire _05402_;
wire _05403_;
wire _05404_;
wire _05405_;
wire _05406_;
wire _05407_;
wire _05408_;
wire _05409_;
wire _05410_;
wire _05411_;
wire _05412_;
wire _05413_;
wire _05414_;
wire _05415_;
wire _05416_;
wire _05417_;
wire _05418_;
wire _05419_;
wire _05420_;
wire _05421_;
wire _05422_;
wire _05423_;
wire _05424_;
wire _05425_;
wire _05426_;
wire _05427_;
wire _05428_;
wire _05429_;
wire _05430_;
wire _05431_;
wire _05432_;
wire _05433_;
wire _05434_;
wire _05435_;
wire _05436_;
wire _05437_;
wire _05438_;
wire _05439_;
wire _05440_;
wire _05441_;
wire _05442_;
wire _05443_;
wire _05444_;
wire _05445_;
wire _05446_;
wire _05447_;
wire _05448_;
wire _05449_;
wire _05450_;
wire _05451_;
wire _05452_;
wire _05453_;
wire _05454_;
wire _05455_;
wire _05456_;
wire _05457_;
wire _05458_;
wire _05459_;
wire _05460_;
wire _05461_;
wire _05462_;
wire _05463_;
wire _05464_;
wire _05465_;
wire _05466_;
wire _05467_;
wire _05468_;
wire _05469_;
wire _05470_;
wire _05471_;
wire _05472_;
wire _05473_;
wire _05474_;
wire _05475_;
wire _05476_;
wire _05477_;
wire _05478_;
wire _05479_;
wire _05480_;
wire _05481_;
wire _05482_;
wire _05483_;
wire _05484_;
wire _05485_;
wire _05486_;
wire _05487_;
wire _05488_;
wire _05489_;
wire _05490_;
wire _05491_;
wire _05492_;
wire _05493_;
wire _05494_;
wire _05495_;
wire _05496_;
wire _05497_;
wire _05498_;
wire _05499_;
wire _05500_;
wire _05501_;
wire _05502_;
wire _05503_;
wire _05504_;
wire _05505_;
wire _05506_;
wire _05507_;
wire _05508_;
wire _05509_;
wire _05510_;
wire _05511_;
wire _05512_;
wire _05513_;
wire _05514_;
wire _05515_;
wire _05516_;
wire _05517_;
wire _05518_;
wire _05519_;
wire _05520_;
wire _05521_;
wire _05522_;
wire _05523_;
wire _05524_;
wire _05525_;
wire _05526_;
wire _05527_;
wire _05528_;
wire _05529_;
wire _05530_;
wire _05531_;
wire _05532_;
wire _05533_;
wire _05534_;
wire _05535_;
wire _05536_;
wire _05537_;
wire _05538_;
wire _05539_;
wire _05540_;
wire _05541_;
wire _05542_;
wire _05543_;
wire _05544_;
wire _05545_;
wire _05546_;
wire _05547_;
wire _05548_;
wire _05549_;
wire _05550_;
wire _05551_;
wire _05552_;
wire _05553_;
wire _05554_;
wire _05555_;
wire _05556_;
wire _05557_;
wire _05558_;
wire _05559_;
wire _05560_;
wire _05561_;
wire _05562_;
wire _05563_;
wire _05564_;
wire _05565_;
wire _05566_;
wire _05567_;
wire _05568_;
wire _05569_;
wire _05570_;
wire _05571_;
wire _05572_;
wire _05573_;
wire _05574_;
wire _05575_;
wire _05576_;
wire _05577_;
wire _05578_;
wire _05579_;
wire _05580_;
wire _05581_;
wire _05582_;
wire _05583_;
wire _05584_;
wire _05585_;
wire _05586_;
wire _05587_;
wire _05588_;
wire _05589_;
wire _05590_;
wire _05591_;
wire _05592_;
wire _05593_;
wire _05594_;
wire _05595_;
wire _05596_;
wire _05597_;
wire _05598_;
wire _05599_;
wire _05600_;
wire _05601_;
wire _05602_;
wire _05603_;
wire _05604_;
wire _05605_;
wire _05606_;
wire _05607_;
wire _05608_;
wire _05609_;
wire _05610_;
wire _05611_;
wire _05612_;
wire _05613_;
wire _05614_;
wire _05615_;
wire _05616_;
wire _05617_;
wire _05618_;
wire _05619_;
wire _05620_;
wire _05621_;
wire _05622_;
wire _05623_;
wire _05624_;
wire _05625_;
wire _05626_;
wire _05627_;
wire _05628_;
wire _05629_;
wire _05630_;
wire _05631_;
wire _05632_;
wire _05633_;
wire _05634_;
wire _05635_;
wire _05636_;
wire _05637_;
wire _05638_;
wire _05639_;
wire _05640_;
wire _05641_;
wire _05642_;
wire _05643_;
wire _05644_;
wire _05645_;
wire _05646_;
wire _05647_;
wire _05648_;
wire _05649_;
wire _05650_;
wire _05651_;
wire _05652_;
wire _05653_;
wire _05654_;
wire _05655_;
wire _05656_;
wire _05657_;
wire _05658_;
wire _05659_;
wire _05660_;
wire _05661_;
wire _05662_;
wire _05663_;
wire _05664_;
wire _05665_;
wire _05666_;
wire _05667_;
wire _05668_;
wire _05669_;
wire _05670_;
wire _05671_;
wire _05672_;
wire _05673_;
wire _05674_;
wire _05675_;
wire _05676_;
wire _05677_;
wire _05678_;
wire _05679_;
wire _05680_;
wire _05681_;
wire _05682_;
wire _05683_;
wire \sresult[0][0] ;
wire \sresult[0][10] ;
wire \sresult[0][11] ;
wire \sresult[0][1] ;
wire \sresult[0][2] ;
wire \sresult[0][3] ;
wire \sresult[0][4] ;
wire \sresult[0][5] ;
wire \sresult[0][6] ;
wire \sresult[0][7] ;
wire \sresult[0][8] ;
wire \sresult[0][9] ;
wire \sresult[10][0] ;
wire \sresult[10][10] ;
wire \sresult[10][11] ;
wire \sresult[10][1] ;
wire \sresult[10][2] ;
wire \sresult[10][3] ;
wire \sresult[10][4] ;
wire \sresult[10][5] ;
wire \sresult[10][6] ;
wire \sresult[10][7] ;
wire \sresult[10][8] ;
wire \sresult[10][9] ;
wire \sresult[11][0] ;
wire \sresult[11][10] ;
wire \sresult[11][11] ;
wire \sresult[11][1] ;
wire \sresult[11][2] ;
wire \sresult[11][3] ;
wire \sresult[11][4] ;
wire \sresult[11][5] ;
wire \sresult[11][6] ;
wire \sresult[11][7] ;
wire \sresult[11][8] ;
wire \sresult[11][9] ;
wire \sresult[12][0] ;
wire \sresult[12][10] ;
wire \sresult[12][11] ;
wire \sresult[12][1] ;
wire \sresult[12][2] ;
wire \sresult[12][3] ;
wire \sresult[12][4] ;
wire \sresult[12][5] ;
wire \sresult[12][6] ;
wire \sresult[12][7] ;
wire \sresult[12][8] ;
wire \sresult[12][9] ;
wire \sresult[13][0] ;
wire \sresult[13][10] ;
wire \sresult[13][11] ;
wire \sresult[13][1] ;
wire \sresult[13][2] ;
wire \sresult[13][3] ;
wire \sresult[13][4] ;
wire \sresult[13][5] ;
wire \sresult[13][6] ;
wire \sresult[13][7] ;
wire \sresult[13][8] ;
wire \sresult[13][9] ;
wire \sresult[14][0] ;
wire \sresult[14][10] ;
wire \sresult[14][11] ;
wire \sresult[14][1] ;
wire \sresult[14][2] ;
wire \sresult[14][3] ;
wire \sresult[14][4] ;
wire \sresult[14][5] ;
wire \sresult[14][6] ;
wire \sresult[14][7] ;
wire \sresult[14][8] ;
wire \sresult[14][9] ;
wire \sresult[15][0] ;
wire \sresult[15][10] ;
wire \sresult[15][11] ;
wire \sresult[15][1] ;
wire \sresult[15][2] ;
wire \sresult[15][3] ;
wire \sresult[15][4] ;
wire \sresult[15][5] ;
wire \sresult[15][6] ;
wire \sresult[15][7] ;
wire \sresult[15][8] ;
wire \sresult[15][9] ;
wire \sresult[16][0] ;
wire \sresult[16][10] ;
wire \sresult[16][11] ;
wire \sresult[16][1] ;
wire \sresult[16][2] ;
wire \sresult[16][3] ;
wire \sresult[16][4] ;
wire \sresult[16][5] ;
wire \sresult[16][6] ;
wire \sresult[16][7] ;
wire \sresult[16][8] ;
wire \sresult[16][9] ;
wire \sresult[17][0] ;
wire \sresult[17][10] ;
wire \sresult[17][11] ;
wire \sresult[17][1] ;
wire \sresult[17][2] ;
wire \sresult[17][3] ;
wire \sresult[17][4] ;
wire \sresult[17][5] ;
wire \sresult[17][6] ;
wire \sresult[17][7] ;
wire \sresult[17][8] ;
wire \sresult[17][9] ;
wire \sresult[18][0] ;
wire \sresult[18][10] ;
wire \sresult[18][11] ;
wire \sresult[18][1] ;
wire \sresult[18][2] ;
wire \sresult[18][3] ;
wire \sresult[18][4] ;
wire \sresult[18][5] ;
wire \sresult[18][6] ;
wire \sresult[18][7] ;
wire \sresult[18][8] ;
wire \sresult[18][9] ;
wire \sresult[19][0] ;
wire \sresult[19][10] ;
wire \sresult[19][11] ;
wire \sresult[19][1] ;
wire \sresult[19][2] ;
wire \sresult[19][3] ;
wire \sresult[19][4] ;
wire \sresult[19][5] ;
wire \sresult[19][6] ;
wire \sresult[19][7] ;
wire \sresult[19][8] ;
wire \sresult[19][9] ;
wire \sresult[1][0] ;
wire \sresult[1][10] ;
wire \sresult[1][11] ;
wire \sresult[1][1] ;
wire \sresult[1][2] ;
wire \sresult[1][3] ;
wire \sresult[1][4] ;
wire \sresult[1][5] ;
wire \sresult[1][6] ;
wire \sresult[1][7] ;
wire \sresult[1][8] ;
wire \sresult[1][9] ;
wire \sresult[20][0] ;
wire \sresult[20][10] ;
wire \sresult[20][11] ;
wire \sresult[20][1] ;
wire \sresult[20][2] ;
wire \sresult[20][3] ;
wire \sresult[20][4] ;
wire \sresult[20][5] ;
wire \sresult[20][6] ;
wire \sresult[20][7] ;
wire \sresult[20][8] ;
wire \sresult[20][9] ;
wire \sresult[21][0] ;
wire \sresult[21][10] ;
wire \sresult[21][11] ;
wire \sresult[21][1] ;
wire \sresult[21][2] ;
wire \sresult[21][3] ;
wire \sresult[21][4] ;
wire \sresult[21][5] ;
wire \sresult[21][6] ;
wire \sresult[21][7] ;
wire \sresult[21][8] ;
wire \sresult[21][9] ;
wire \sresult[22][0] ;
wire \sresult[22][10] ;
wire \sresult[22][11] ;
wire \sresult[22][1] ;
wire \sresult[22][2] ;
wire \sresult[22][3] ;
wire \sresult[22][4] ;
wire \sresult[22][5] ;
wire \sresult[22][6] ;
wire \sresult[22][7] ;
wire \sresult[22][8] ;
wire \sresult[22][9] ;
wire \sresult[23][0] ;
wire \sresult[23][10] ;
wire \sresult[23][11] ;
wire \sresult[23][1] ;
wire \sresult[23][2] ;
wire \sresult[23][3] ;
wire \sresult[23][4] ;
wire \sresult[23][5] ;
wire \sresult[23][6] ;
wire \sresult[23][7] ;
wire \sresult[23][8] ;
wire \sresult[23][9] ;
wire \sresult[24][0] ;
wire \sresult[24][10] ;
wire \sresult[24][11] ;
wire \sresult[24][1] ;
wire \sresult[24][2] ;
wire \sresult[24][3] ;
wire \sresult[24][4] ;
wire \sresult[24][5] ;
wire \sresult[24][6] ;
wire \sresult[24][7] ;
wire \sresult[24][8] ;
wire \sresult[24][9] ;
wire \sresult[25][0] ;
wire \sresult[25][10] ;
wire \sresult[25][11] ;
wire \sresult[25][1] ;
wire \sresult[25][2] ;
wire \sresult[25][3] ;
wire \sresult[25][4] ;
wire \sresult[25][5] ;
wire \sresult[25][6] ;
wire \sresult[25][7] ;
wire \sresult[25][8] ;
wire \sresult[25][9] ;
wire \sresult[26][0] ;
wire \sresult[26][10] ;
wire \sresult[26][11] ;
wire \sresult[26][1] ;
wire \sresult[26][2] ;
wire \sresult[26][3] ;
wire \sresult[26][4] ;
wire \sresult[26][5] ;
wire \sresult[26][6] ;
wire \sresult[26][7] ;
wire \sresult[26][8] ;
wire \sresult[26][9] ;
wire \sresult[27][0] ;
wire \sresult[27][10] ;
wire \sresult[27][11] ;
wire \sresult[27][1] ;
wire \sresult[27][2] ;
wire \sresult[27][3] ;
wire \sresult[27][4] ;
wire \sresult[27][5] ;
wire \sresult[27][6] ;
wire \sresult[27][7] ;
wire \sresult[27][8] ;
wire \sresult[27][9] ;
wire \sresult[28][0] ;
wire \sresult[28][10] ;
wire \sresult[28][11] ;
wire \sresult[28][1] ;
wire \sresult[28][2] ;
wire \sresult[28][3] ;
wire \sresult[28][4] ;
wire \sresult[28][5] ;
wire \sresult[28][6] ;
wire \sresult[28][7] ;
wire \sresult[28][8] ;
wire \sresult[28][9] ;
wire \sresult[29][0] ;
wire \sresult[29][10] ;
wire \sresult[29][11] ;
wire \sresult[29][1] ;
wire \sresult[29][2] ;
wire \sresult[29][3] ;
wire \sresult[29][4] ;
wire \sresult[29][5] ;
wire \sresult[29][6] ;
wire \sresult[29][7] ;
wire \sresult[29][8] ;
wire \sresult[29][9] ;
wire \sresult[2][0] ;
wire \sresult[2][10] ;
wire \sresult[2][11] ;
wire \sresult[2][1] ;
wire \sresult[2][2] ;
wire \sresult[2][3] ;
wire \sresult[2][4] ;
wire \sresult[2][5] ;
wire \sresult[2][6] ;
wire \sresult[2][7] ;
wire \sresult[2][8] ;
wire \sresult[2][9] ;
wire \sresult[30][0] ;
wire \sresult[30][10] ;
wire \sresult[30][11] ;
wire \sresult[30][1] ;
wire \sresult[30][2] ;
wire \sresult[30][3] ;
wire \sresult[30][4] ;
wire \sresult[30][5] ;
wire \sresult[30][6] ;
wire \sresult[30][7] ;
wire \sresult[30][8] ;
wire \sresult[30][9] ;
wire \sresult[31][0] ;
wire \sresult[31][10] ;
wire \sresult[31][11] ;
wire \sresult[31][1] ;
wire \sresult[31][2] ;
wire \sresult[31][3] ;
wire \sresult[31][4] ;
wire \sresult[31][5] ;
wire \sresult[31][6] ;
wire \sresult[31][7] ;
wire \sresult[31][8] ;
wire \sresult[31][9] ;
wire \sresult[32][0] ;
wire \sresult[32][10] ;
wire \sresult[32][11] ;
wire \sresult[32][1] ;
wire \sresult[32][2] ;
wire \sresult[32][3] ;
wire \sresult[32][4] ;
wire \sresult[32][5] ;
wire \sresult[32][6] ;
wire \sresult[32][7] ;
wire \sresult[32][8] ;
wire \sresult[32][9] ;
wire \sresult[33][0] ;
wire \sresult[33][10] ;
wire \sresult[33][11] ;
wire \sresult[33][1] ;
wire \sresult[33][2] ;
wire \sresult[33][3] ;
wire \sresult[33][4] ;
wire \sresult[33][5] ;
wire \sresult[33][6] ;
wire \sresult[33][7] ;
wire \sresult[33][8] ;
wire \sresult[33][9] ;
wire \sresult[34][0] ;
wire \sresult[34][10] ;
wire \sresult[34][11] ;
wire \sresult[34][1] ;
wire \sresult[34][2] ;
wire \sresult[34][3] ;
wire \sresult[34][4] ;
wire \sresult[34][5] ;
wire \sresult[34][6] ;
wire \sresult[34][7] ;
wire \sresult[34][8] ;
wire \sresult[34][9] ;
wire \sresult[35][0] ;
wire \sresult[35][10] ;
wire \sresult[35][11] ;
wire \sresult[35][1] ;
wire \sresult[35][2] ;
wire \sresult[35][3] ;
wire \sresult[35][4] ;
wire \sresult[35][5] ;
wire \sresult[35][6] ;
wire \sresult[35][7] ;
wire \sresult[35][8] ;
wire \sresult[35][9] ;
wire \sresult[36][0] ;
wire \sresult[36][10] ;
wire \sresult[36][11] ;
wire \sresult[36][1] ;
wire \sresult[36][2] ;
wire \sresult[36][3] ;
wire \sresult[36][4] ;
wire \sresult[36][5] ;
wire \sresult[36][6] ;
wire \sresult[36][7] ;
wire \sresult[36][8] ;
wire \sresult[36][9] ;
wire \sresult[37][0] ;
wire \sresult[37][10] ;
wire \sresult[37][11] ;
wire \sresult[37][1] ;
wire \sresult[37][2] ;
wire \sresult[37][3] ;
wire \sresult[37][4] ;
wire \sresult[37][5] ;
wire \sresult[37][6] ;
wire \sresult[37][7] ;
wire \sresult[37][8] ;
wire \sresult[37][9] ;
wire \sresult[38][0] ;
wire \sresult[38][10] ;
wire \sresult[38][11] ;
wire \sresult[38][1] ;
wire \sresult[38][2] ;
wire \sresult[38][3] ;
wire \sresult[38][4] ;
wire \sresult[38][5] ;
wire \sresult[38][6] ;
wire \sresult[38][7] ;
wire \sresult[38][8] ;
wire \sresult[38][9] ;
wire \sresult[39][0] ;
wire \sresult[39][10] ;
wire \sresult[39][11] ;
wire \sresult[39][1] ;
wire \sresult[39][2] ;
wire \sresult[39][3] ;
wire \sresult[39][4] ;
wire \sresult[39][5] ;
wire \sresult[39][6] ;
wire \sresult[39][7] ;
wire \sresult[39][8] ;
wire \sresult[39][9] ;
wire \sresult[3][0] ;
wire \sresult[3][10] ;
wire \sresult[3][11] ;
wire \sresult[3][1] ;
wire \sresult[3][2] ;
wire \sresult[3][3] ;
wire \sresult[3][4] ;
wire \sresult[3][5] ;
wire \sresult[3][6] ;
wire \sresult[3][7] ;
wire \sresult[3][8] ;
wire \sresult[3][9] ;
wire \sresult[40][0] ;
wire \sresult[40][10] ;
wire \sresult[40][11] ;
wire \sresult[40][1] ;
wire \sresult[40][2] ;
wire \sresult[40][3] ;
wire \sresult[40][4] ;
wire \sresult[40][5] ;
wire \sresult[40][6] ;
wire \sresult[40][7] ;
wire \sresult[40][8] ;
wire \sresult[40][9] ;
wire \sresult[41][0] ;
wire \sresult[41][10] ;
wire \sresult[41][11] ;
wire \sresult[41][1] ;
wire \sresult[41][2] ;
wire \sresult[41][3] ;
wire \sresult[41][4] ;
wire \sresult[41][5] ;
wire \sresult[41][6] ;
wire \sresult[41][7] ;
wire \sresult[41][8] ;
wire \sresult[41][9] ;
wire \sresult[42][0] ;
wire \sresult[42][10] ;
wire \sresult[42][11] ;
wire \sresult[42][1] ;
wire \sresult[42][2] ;
wire \sresult[42][3] ;
wire \sresult[42][4] ;
wire \sresult[42][5] ;
wire \sresult[42][6] ;
wire \sresult[42][7] ;
wire \sresult[42][8] ;
wire \sresult[42][9] ;
wire \sresult[43][0] ;
wire \sresult[43][10] ;
wire \sresult[43][11] ;
wire \sresult[43][1] ;
wire \sresult[43][2] ;
wire \sresult[43][3] ;
wire \sresult[43][4] ;
wire \sresult[43][5] ;
wire \sresult[43][6] ;
wire \sresult[43][7] ;
wire \sresult[43][8] ;
wire \sresult[43][9] ;
wire \sresult[44][0] ;
wire \sresult[44][10] ;
wire \sresult[44][11] ;
wire \sresult[44][1] ;
wire \sresult[44][2] ;
wire \sresult[44][3] ;
wire \sresult[44][4] ;
wire \sresult[44][5] ;
wire \sresult[44][6] ;
wire \sresult[44][7] ;
wire \sresult[44][8] ;
wire \sresult[44][9] ;
wire \sresult[45][0] ;
wire \sresult[45][10] ;
wire \sresult[45][11] ;
wire \sresult[45][1] ;
wire \sresult[45][2] ;
wire \sresult[45][3] ;
wire \sresult[45][4] ;
wire \sresult[45][5] ;
wire \sresult[45][6] ;
wire \sresult[45][7] ;
wire \sresult[45][8] ;
wire \sresult[45][9] ;
wire \sresult[46][0] ;
wire \sresult[46][10] ;
wire \sresult[46][11] ;
wire \sresult[46][1] ;
wire \sresult[46][2] ;
wire \sresult[46][3] ;
wire \sresult[46][4] ;
wire \sresult[46][5] ;
wire \sresult[46][6] ;
wire \sresult[46][7] ;
wire \sresult[46][8] ;
wire \sresult[46][9] ;
wire \sresult[47][0] ;
wire \sresult[47][10] ;
wire \sresult[47][11] ;
wire \sresult[47][1] ;
wire \sresult[47][2] ;
wire \sresult[47][3] ;
wire \sresult[47][4] ;
wire \sresult[47][5] ;
wire \sresult[47][6] ;
wire \sresult[47][7] ;
wire \sresult[47][8] ;
wire \sresult[47][9] ;
wire \sresult[48][0] ;
wire \sresult[48][10] ;
wire \sresult[48][11] ;
wire \sresult[48][1] ;
wire \sresult[48][2] ;
wire \sresult[48][3] ;
wire \sresult[48][4] ;
wire \sresult[48][5] ;
wire \sresult[48][6] ;
wire \sresult[48][7] ;
wire \sresult[48][8] ;
wire \sresult[48][9] ;
wire \sresult[49][0] ;
wire \sresult[49][10] ;
wire \sresult[49][11] ;
wire \sresult[49][1] ;
wire \sresult[49][2] ;
wire \sresult[49][3] ;
wire \sresult[49][4] ;
wire \sresult[49][5] ;
wire \sresult[49][6] ;
wire \sresult[49][7] ;
wire \sresult[49][8] ;
wire \sresult[49][9] ;
wire \sresult[4][0] ;
wire \sresult[4][10] ;
wire \sresult[4][11] ;
wire \sresult[4][1] ;
wire \sresult[4][2] ;
wire \sresult[4][3] ;
wire \sresult[4][4] ;
wire \sresult[4][5] ;
wire \sresult[4][6] ;
wire \sresult[4][7] ;
wire \sresult[4][8] ;
wire \sresult[4][9] ;
wire \sresult[50][0] ;
wire \sresult[50][10] ;
wire \sresult[50][11] ;
wire \sresult[50][1] ;
wire \sresult[50][2] ;
wire \sresult[50][3] ;
wire \sresult[50][4] ;
wire \sresult[50][5] ;
wire \sresult[50][6] ;
wire \sresult[50][7] ;
wire \sresult[50][8] ;
wire \sresult[50][9] ;
wire \sresult[51][0] ;
wire \sresult[51][10] ;
wire \sresult[51][11] ;
wire \sresult[51][1] ;
wire \sresult[51][2] ;
wire \sresult[51][3] ;
wire \sresult[51][4] ;
wire \sresult[51][5] ;
wire \sresult[51][6] ;
wire \sresult[51][7] ;
wire \sresult[51][8] ;
wire \sresult[51][9] ;
wire \sresult[52][0] ;
wire \sresult[52][10] ;
wire \sresult[52][11] ;
wire \sresult[52][1] ;
wire \sresult[52][2] ;
wire \sresult[52][3] ;
wire \sresult[52][4] ;
wire \sresult[52][5] ;
wire \sresult[52][6] ;
wire \sresult[52][7] ;
wire \sresult[52][8] ;
wire \sresult[52][9] ;
wire \sresult[53][0] ;
wire \sresult[53][10] ;
wire \sresult[53][11] ;
wire \sresult[53][1] ;
wire \sresult[53][2] ;
wire \sresult[53][3] ;
wire \sresult[53][4] ;
wire \sresult[53][5] ;
wire \sresult[53][6] ;
wire \sresult[53][7] ;
wire \sresult[53][8] ;
wire \sresult[53][9] ;
wire \sresult[54][0] ;
wire \sresult[54][10] ;
wire \sresult[54][11] ;
wire \sresult[54][1] ;
wire \sresult[54][2] ;
wire \sresult[54][3] ;
wire \sresult[54][4] ;
wire \sresult[54][5] ;
wire \sresult[54][6] ;
wire \sresult[54][7] ;
wire \sresult[54][8] ;
wire \sresult[54][9] ;
wire \sresult[55][0] ;
wire \sresult[55][10] ;
wire \sresult[55][11] ;
wire \sresult[55][1] ;
wire \sresult[55][2] ;
wire \sresult[55][3] ;
wire \sresult[55][4] ;
wire \sresult[55][5] ;
wire \sresult[55][6] ;
wire \sresult[55][7] ;
wire \sresult[55][8] ;
wire \sresult[55][9] ;
wire \sresult[56][0] ;
wire \sresult[56][10] ;
wire \sresult[56][11] ;
wire \sresult[56][1] ;
wire \sresult[56][2] ;
wire \sresult[56][3] ;
wire \sresult[56][4] ;
wire \sresult[56][5] ;
wire \sresult[56][6] ;
wire \sresult[56][7] ;
wire \sresult[56][8] ;
wire \sresult[56][9] ;
wire \sresult[57][0] ;
wire \sresult[57][10] ;
wire \sresult[57][11] ;
wire \sresult[57][1] ;
wire \sresult[57][2] ;
wire \sresult[57][3] ;
wire \sresult[57][4] ;
wire \sresult[57][5] ;
wire \sresult[57][6] ;
wire \sresult[57][7] ;
wire \sresult[57][8] ;
wire \sresult[57][9] ;
wire \sresult[58][0] ;
wire \sresult[58][10] ;
wire \sresult[58][11] ;
wire \sresult[58][1] ;
wire \sresult[58][2] ;
wire \sresult[58][3] ;
wire \sresult[58][4] ;
wire \sresult[58][5] ;
wire \sresult[58][6] ;
wire \sresult[58][7] ;
wire \sresult[58][8] ;
wire \sresult[58][9] ;
wire \sresult[59][0] ;
wire \sresult[59][10] ;
wire \sresult[59][11] ;
wire \sresult[59][1] ;
wire \sresult[59][2] ;
wire \sresult[59][3] ;
wire \sresult[59][4] ;
wire \sresult[59][5] ;
wire \sresult[59][6] ;
wire \sresult[59][7] ;
wire \sresult[59][8] ;
wire \sresult[59][9] ;
wire \sresult[5][0] ;
wire \sresult[5][10] ;
wire \sresult[5][11] ;
wire \sresult[5][1] ;
wire \sresult[5][2] ;
wire \sresult[5][3] ;
wire \sresult[5][4] ;
wire \sresult[5][5] ;
wire \sresult[5][6] ;
wire \sresult[5][7] ;
wire \sresult[5][8] ;
wire \sresult[5][9] ;
wire \sresult[60][0] ;
wire \sresult[60][10] ;
wire \sresult[60][11] ;
wire \sresult[60][1] ;
wire \sresult[60][2] ;
wire \sresult[60][3] ;
wire \sresult[60][4] ;
wire \sresult[60][5] ;
wire \sresult[60][6] ;
wire \sresult[60][7] ;
wire \sresult[60][8] ;
wire \sresult[60][9] ;
wire \sresult[61][0] ;
wire \sresult[61][10] ;
wire \sresult[61][11] ;
wire \sresult[61][1] ;
wire \sresult[61][2] ;
wire \sresult[61][3] ;
wire \sresult[61][4] ;
wire \sresult[61][5] ;
wire \sresult[61][6] ;
wire \sresult[61][7] ;
wire \sresult[61][8] ;
wire \sresult[61][9] ;
wire \sresult[62][0] ;
wire \sresult[62][10] ;
wire \sresult[62][11] ;
wire \sresult[62][1] ;
wire \sresult[62][2] ;
wire \sresult[62][3] ;
wire \sresult[62][4] ;
wire \sresult[62][5] ;
wire \sresult[62][6] ;
wire \sresult[62][7] ;
wire \sresult[62][8] ;
wire \sresult[62][9] ;
wire \sresult[6][0] ;
wire \sresult[6][10] ;
wire \sresult[6][11] ;
wire \sresult[6][1] ;
wire \sresult[6][2] ;
wire \sresult[6][3] ;
wire \sresult[6][4] ;
wire \sresult[6][5] ;
wire \sresult[6][6] ;
wire \sresult[6][7] ;
wire \sresult[6][8] ;
wire \sresult[6][9] ;
wire \sresult[7][0] ;
wire \sresult[7][10] ;
wire \sresult[7][11] ;
wire \sresult[7][1] ;
wire \sresult[7][2] ;
wire \sresult[7][3] ;
wire \sresult[7][4] ;
wire \sresult[7][5] ;
wire \sresult[7][6] ;
wire \sresult[7][7] ;
wire \sresult[7][8] ;
wire \sresult[7][9] ;
wire \sresult[8][0] ;
wire \sresult[8][10] ;
wire \sresult[8][11] ;
wire \sresult[8][1] ;
wire \sresult[8][2] ;
wire \sresult[8][3] ;
wire \sresult[8][4] ;
wire \sresult[8][5] ;
wire \sresult[8][6] ;
wire \sresult[8][7] ;
wire \sresult[8][8] ;
wire \sresult[8][9] ;
wire \sresult[9][0] ;
wire \sresult[9][10] ;
wire \sresult[9][11] ;
wire \sresult[9][1] ;
wire \sresult[9][2] ;
wire \sresult[9][3] ;
wire \sresult[9][4] ;
wire \sresult[9][5] ;
wire \sresult[9][6] ;
wire \sresult[9][7] ;
wire \sresult[9][8] ;
wire \sresult[9][9] ;

BUF_X4 _05684_ (
  .A(douten),
  .Z(_00769_)
);

BUF_X16 _05685_ (
  .A(_00769_),
  .Z(_00770_)
);

BUF_X4 _05686_ (
  .A(ena),
  .Z(_00771_)
);

NAND2_X2 _05687_ (
  .A1(_00770_),
  .A2(_00771_),
  .ZN(_00772_)
);

NAND2_X1 _05688_ (
  .A1(_00772_),
  .A2(\sresult[0][0] ),
  .ZN(_00773_)
);

INV_X1 _05689_ (
  .A(din_77[0]),
  .ZN(_00774_)
);

BUF_X2 _05690_ (
  .A(_00772_),
  .Z(_00775_)
);

OAI21_X1 _05691_ (
  .A(_00773_),
  .B1(_00774_),
  .B2(_00775_),
  .ZN(_00000_)
);

NAND2_X1 _05692_ (
  .A1(_00772_),
  .A2(\sresult[0][1] ),
  .ZN(_00776_)
);

INV_X1 _05693_ (
  .A(din_77[1]),
  .ZN(_00777_)
);

OAI21_X1 _05694_ (
  .A(_00776_),
  .B1(_00777_),
  .B2(_00775_),
  .ZN(_00001_)
);

BUF_X2 _05695_ (
  .A(_00772_),
  .Z(_00778_)
);

NAND2_X1 _05696_ (
  .A1(_00778_),
  .A2(\sresult[0][2] ),
  .ZN(_00779_)
);

INV_X1 _05697_ (
  .A(din_77[2]),
  .ZN(_00780_)
);

OAI21_X1 _05698_ (
  .A(_00779_),
  .B1(_00780_),
  .B2(_00775_),
  .ZN(_00002_)
);

NAND2_X1 _05699_ (
  .A1(_00772_),
  .A2(\sresult[0][3] ),
  .ZN(_00781_)
);

INV_X1 _05700_ (
  .A(din_77[3]),
  .ZN(_00782_)
);

OAI21_X1 _05701_ (
  .A(_00781_),
  .B1(_00782_),
  .B2(_00775_),
  .ZN(_00003_)
);

NAND2_X1 _05702_ (
  .A1(_00778_),
  .A2(\sresult[0][4] ),
  .ZN(_00783_)
);

INV_X1 _05703_ (
  .A(din_77[4]),
  .ZN(_00784_)
);

OAI21_X1 _05704_ (
  .A(_00783_),
  .B1(_00784_),
  .B2(_00775_),
  .ZN(_00004_)
);

NAND2_X1 _05705_ (
  .A1(_00778_),
  .A2(\sresult[0][5] ),
  .ZN(_00785_)
);

INV_X1 _05706_ (
  .A(din_77[5]),
  .ZN(_00786_)
);

OAI21_X1 _05707_ (
  .A(_00785_),
  .B1(_00786_),
  .B2(_00778_),
  .ZN(_00005_)
);

NAND2_X1 _05708_ (
  .A1(_00778_),
  .A2(\sresult[0][6] ),
  .ZN(_00787_)
);

INV_X1 _05709_ (
  .A(din_77[6]),
  .ZN(_00788_)
);

OAI21_X1 _05710_ (
  .A(_00787_),
  .B1(_00788_),
  .B2(_00775_),
  .ZN(_00006_)
);

NAND2_X1 _05711_ (
  .A1(_00778_),
  .A2(\sresult[0][7] ),
  .ZN(_00789_)
);

INV_X1 _05712_ (
  .A(din_77[7]),
  .ZN(_00790_)
);

OAI21_X1 _05713_ (
  .A(_00789_),
  .B1(_00790_),
  .B2(_00775_),
  .ZN(_00007_)
);

NAND2_X1 _05714_ (
  .A1(_00778_),
  .A2(\sresult[0][8] ),
  .ZN(_00791_)
);

INV_X1 _05715_ (
  .A(din_77[8]),
  .ZN(_00792_)
);

OAI21_X1 _05716_ (
  .A(_00791_),
  .B1(_00792_),
  .B2(_00775_),
  .ZN(_00008_)
);

NAND2_X1 _05717_ (
  .A1(_00778_),
  .A2(\sresult[0][9] ),
  .ZN(_00793_)
);

INV_X1 _05718_ (
  .A(din_77[9]),
  .ZN(_00794_)
);

OAI21_X1 _05719_ (
  .A(_00793_),
  .B1(_00794_),
  .B2(_00775_),
  .ZN(_00009_)
);

NAND2_X1 _05720_ (
  .A1(_00772_),
  .A2(\sresult[0][10] ),
  .ZN(_00795_)
);

INV_X1 _05721_ (
  .A(din_77[10]),
  .ZN(_00796_)
);

OAI21_X1 _05722_ (
  .A(_00795_),
  .B1(_00796_),
  .B2(_00778_),
  .ZN(_00010_)
);

NAND2_X1 _05723_ (
  .A1(_00778_),
  .A2(\sresult[0][11] ),
  .ZN(_00797_)
);

INV_X1 _05724_ (
  .A(din_77[11]),
  .ZN(_00798_)
);

OAI21_X1 _05725_ (
  .A(_00797_),
  .B1(_00798_),
  .B2(_00775_),
  .ZN(_00011_)
);

INV_X8 _05726_ (
  .A(_00769_),
  .ZN(_00799_)
);

BUF_X8 _05727_ (
  .A(_00799_),
  .Z(_00800_)
);

BUF_X4 _05728_ (
  .A(_00800_),
  .Z(_00801_)
);

NAND2_X1 _05729_ (
  .A1(_00801_),
  .A2(\sresult[0][0] ),
  .ZN(_00802_)
);

BUF_X8 _05730_ (
  .A(_00770_),
  .Z(_00803_)
);

BUF_X4 _05731_ (
  .A(_00803_),
  .Z(_00804_)
);

NAND2_X1 _05732_ (
  .A1(_00804_),
  .A2(din_76[0]),
  .ZN(_00805_)
);

NAND2_X1 _05733_ (
  .A1(_00802_),
  .A2(_00805_),
  .ZN(_00806_)
);

BUF_X2 _05734_ (
  .A(_00771_),
  .Z(_00807_)
);

BUF_X2 _05735_ (
  .A(_00807_),
  .Z(_00808_)
);

NAND2_X1 _05736_ (
  .A1(_00806_),
  .A2(_00808_),
  .ZN(_00809_)
);

INV_X8 _05737_ (
  .A(_00771_),
  .ZN(_00810_)
);

BUF_X8 _05738_ (
  .A(_00810_),
  .Z(_00811_)
);

CLKBUF_X2 _05739_ (
  .A(_00811_),
  .Z(_00812_)
);

NAND2_X1 _05740_ (
  .A1(_00812_),
  .A2(\sresult[1][0] ),
  .ZN(_00813_)
);

NAND2_X1 _05741_ (
  .A1(_00809_),
  .A2(_00813_),
  .ZN(_00012_)
);

BUF_X4 _05742_ (
  .A(_00799_),
  .Z(_00814_)
);

BUF_X4 _05743_ (
  .A(_00814_),
  .Z(_00815_)
);

NAND2_X1 _05744_ (
  .A1(_00815_),
  .A2(\sresult[0][1] ),
  .ZN(_00816_)
);

NAND2_X1 _05745_ (
  .A1(_00804_),
  .A2(din_76[1]),
  .ZN(_00817_)
);

NAND2_X1 _05746_ (
  .A1(_00816_),
  .A2(_00817_),
  .ZN(_00818_)
);

NAND2_X1 _05747_ (
  .A1(_00818_),
  .A2(_00808_),
  .ZN(_00819_)
);

BUF_X4 _05748_ (
  .A(_00810_),
  .Z(_00820_)
);

BUF_X2 _05749_ (
  .A(_00820_),
  .Z(_00821_)
);

NAND2_X1 _05750_ (
  .A1(_00821_),
  .A2(\sresult[1][1] ),
  .ZN(_00822_)
);

NAND2_X1 _05751_ (
  .A1(_00819_),
  .A2(_00822_),
  .ZN(_00013_)
);

NAND2_X1 _05752_ (
  .A1(_00815_),
  .A2(\sresult[0][2] ),
  .ZN(_00823_)
);

NAND2_X1 _05753_ (
  .A1(_00804_),
  .A2(din_76[2]),
  .ZN(_00824_)
);

NAND2_X1 _05754_ (
  .A1(_00823_),
  .A2(_00824_),
  .ZN(_00825_)
);

NAND2_X1 _05755_ (
  .A1(_00825_),
  .A2(_00808_),
  .ZN(_00826_)
);

NAND2_X1 _05756_ (
  .A1(_00821_),
  .A2(\sresult[1][2] ),
  .ZN(_00827_)
);

NAND2_X1 _05757_ (
  .A1(_00826_),
  .A2(_00827_),
  .ZN(_00014_)
);

NAND2_X1 _05758_ (
  .A1(_00815_),
  .A2(\sresult[0][3] ),
  .ZN(_00828_)
);

NAND2_X1 _05759_ (
  .A1(_00804_),
  .A2(din_76[3]),
  .ZN(_00829_)
);

NAND2_X1 _05760_ (
  .A1(_00828_),
  .A2(_00829_),
  .ZN(_00830_)
);

NAND2_X1 _05761_ (
  .A1(_00830_),
  .A2(_00808_),
  .ZN(_00831_)
);

NAND2_X1 _05762_ (
  .A1(_00821_),
  .A2(\sresult[1][3] ),
  .ZN(_00832_)
);

NAND2_X1 _05763_ (
  .A1(_00831_),
  .A2(_00832_),
  .ZN(_00015_)
);

NAND2_X1 _05764_ (
  .A1(_00815_),
  .A2(\sresult[0][4] ),
  .ZN(_00833_)
);

NAND2_X1 _05765_ (
  .A1(_00804_),
  .A2(din_76[4]),
  .ZN(_00834_)
);

NAND2_X1 _05766_ (
  .A1(_00833_),
  .A2(_00834_),
  .ZN(_00835_)
);

NAND2_X1 _05767_ (
  .A1(_00835_),
  .A2(_00808_),
  .ZN(_00836_)
);

NAND2_X1 _05768_ (
  .A1(_00821_),
  .A2(\sresult[1][4] ),
  .ZN(_00837_)
);

NAND2_X1 _05769_ (
  .A1(_00836_),
  .A2(_00837_),
  .ZN(_00016_)
);

NAND2_X1 _05770_ (
  .A1(_00815_),
  .A2(\sresult[0][5] ),
  .ZN(_00838_)
);

NAND2_X1 _05771_ (
  .A1(_00804_),
  .A2(din_76[5]),
  .ZN(_00839_)
);

NAND2_X1 _05772_ (
  .A1(_00838_),
  .A2(_00839_),
  .ZN(_00840_)
);

NAND2_X1 _05773_ (
  .A1(_00840_),
  .A2(_00808_),
  .ZN(_00841_)
);

NAND2_X1 _05774_ (
  .A1(_00821_),
  .A2(\sresult[1][5] ),
  .ZN(_00842_)
);

NAND2_X1 _05775_ (
  .A1(_00841_),
  .A2(_00842_),
  .ZN(_00017_)
);

NAND2_X1 _05776_ (
  .A1(_00815_),
  .A2(\sresult[0][6] ),
  .ZN(_00843_)
);

NAND2_X1 _05777_ (
  .A1(_00804_),
  .A2(din_76[6]),
  .ZN(_00844_)
);

NAND2_X1 _05778_ (
  .A1(_00843_),
  .A2(_00844_),
  .ZN(_00845_)
);

NAND2_X1 _05779_ (
  .A1(_00845_),
  .A2(_00808_),
  .ZN(_00846_)
);

NAND2_X1 _05780_ (
  .A1(_00821_),
  .A2(\sresult[1][6] ),
  .ZN(_00847_)
);

NAND2_X1 _05781_ (
  .A1(_00846_),
  .A2(_00847_),
  .ZN(_00018_)
);

NAND2_X1 _05782_ (
  .A1(_00815_),
  .A2(\sresult[0][7] ),
  .ZN(_00848_)
);

NAND2_X1 _05783_ (
  .A1(_00804_),
  .A2(din_76[7]),
  .ZN(_00849_)
);

NAND2_X1 _05784_ (
  .A1(_00848_),
  .A2(_00849_),
  .ZN(_00850_)
);

NAND2_X1 _05785_ (
  .A1(_00850_),
  .A2(_00808_),
  .ZN(_00851_)
);

NAND2_X1 _05786_ (
  .A1(_00821_),
  .A2(\sresult[1][7] ),
  .ZN(_00852_)
);

NAND2_X1 _05787_ (
  .A1(_00851_),
  .A2(_00852_),
  .ZN(_00019_)
);

NAND2_X1 _05788_ (
  .A1(_00815_),
  .A2(\sresult[0][8] ),
  .ZN(_00853_)
);

BUF_X4 _05789_ (
  .A(_00803_),
  .Z(_00854_)
);

NAND2_X1 _05790_ (
  .A1(_00854_),
  .A2(din_76[8]),
  .ZN(_00855_)
);

NAND2_X1 _05791_ (
  .A1(_00853_),
  .A2(_00855_),
  .ZN(_00856_)
);

BUF_X2 _05792_ (
  .A(_00807_),
  .Z(_00857_)
);

NAND2_X1 _05793_ (
  .A1(_00856_),
  .A2(_00857_),
  .ZN(_00858_)
);

NAND2_X1 _05794_ (
  .A1(_00821_),
  .A2(\sresult[1][8] ),
  .ZN(_00859_)
);

NAND2_X1 _05795_ (
  .A1(_00858_),
  .A2(_00859_),
  .ZN(_00020_)
);

NAND2_X1 _05796_ (
  .A1(_00815_),
  .A2(\sresult[0][9] ),
  .ZN(_00860_)
);

NAND2_X1 _05797_ (
  .A1(_00854_),
  .A2(din_76[9]),
  .ZN(_00861_)
);

NAND2_X1 _05798_ (
  .A1(_00860_),
  .A2(_00861_),
  .ZN(_00862_)
);

NAND2_X1 _05799_ (
  .A1(_00862_),
  .A2(_00857_),
  .ZN(_00863_)
);

NAND2_X1 _05800_ (
  .A1(_00821_),
  .A2(\sresult[1][9] ),
  .ZN(_00864_)
);

NAND2_X1 _05801_ (
  .A1(_00863_),
  .A2(_00864_),
  .ZN(_00021_)
);

BUF_X4 _05802_ (
  .A(_00814_),
  .Z(_00865_)
);

NAND2_X1 _05803_ (
  .A1(_00865_),
  .A2(\sresult[0][10] ),
  .ZN(_00866_)
);

NAND2_X1 _05804_ (
  .A1(_00854_),
  .A2(din_76[10]),
  .ZN(_00867_)
);

NAND2_X1 _05805_ (
  .A1(_00866_),
  .A2(_00867_),
  .ZN(_00868_)
);

NAND2_X1 _05806_ (
  .A1(_00868_),
  .A2(_00857_),
  .ZN(_00869_)
);

CLKBUF_X2 _05807_ (
  .A(_00820_),
  .Z(_00870_)
);

NAND2_X1 _05808_ (
  .A1(_00870_),
  .A2(\sresult[1][10] ),
  .ZN(_00871_)
);

NAND2_X1 _05809_ (
  .A1(_00869_),
  .A2(_00871_),
  .ZN(_00022_)
);

NAND2_X1 _05810_ (
  .A1(_00865_),
  .A2(\sresult[0][11] ),
  .ZN(_00872_)
);

NAND2_X1 _05811_ (
  .A1(_00854_),
  .A2(din_76[11]),
  .ZN(_00873_)
);

NAND2_X1 _05812_ (
  .A1(_00872_),
  .A2(_00873_),
  .ZN(_00874_)
);

NAND2_X1 _05813_ (
  .A1(_00874_),
  .A2(_00857_),
  .ZN(_00875_)
);

NAND2_X1 _05814_ (
  .A1(_00870_),
  .A2(\sresult[1][11] ),
  .ZN(_00876_)
);

NAND2_X1 _05815_ (
  .A1(_00875_),
  .A2(_00876_),
  .ZN(_00023_)
);

NAND2_X1 _05816_ (
  .A1(_00865_),
  .A2(\sresult[1][0] ),
  .ZN(_00877_)
);

NAND2_X1 _05817_ (
  .A1(_00854_),
  .A2(din_67[0]),
  .ZN(_00878_)
);

NAND2_X1 _05818_ (
  .A1(_00877_),
  .A2(_00878_),
  .ZN(_00879_)
);

NAND2_X1 _05819_ (
  .A1(_00879_),
  .A2(_00857_),
  .ZN(_00880_)
);

NAND2_X1 _05820_ (
  .A1(_00870_),
  .A2(\sresult[2][0] ),
  .ZN(_00881_)
);

NAND2_X1 _05821_ (
  .A1(_00880_),
  .A2(_00881_),
  .ZN(_00024_)
);

NAND2_X1 _05822_ (
  .A1(_00865_),
  .A2(\sresult[1][1] ),
  .ZN(_00882_)
);

NAND2_X1 _05823_ (
  .A1(_00854_),
  .A2(din_67[1]),
  .ZN(_00883_)
);

NAND2_X1 _05824_ (
  .A1(_00882_),
  .A2(_00883_),
  .ZN(_00884_)
);

NAND2_X1 _05825_ (
  .A1(_00884_),
  .A2(_00857_),
  .ZN(_00885_)
);

NAND2_X1 _05826_ (
  .A1(_00870_),
  .A2(\sresult[2][1] ),
  .ZN(_00886_)
);

NAND2_X1 _05827_ (
  .A1(_00885_),
  .A2(_00886_),
  .ZN(_00025_)
);

NAND2_X1 _05828_ (
  .A1(_00865_),
  .A2(\sresult[1][2] ),
  .ZN(_00887_)
);

NAND2_X1 _05829_ (
  .A1(_00854_),
  .A2(din_67[2]),
  .ZN(_00888_)
);

NAND2_X1 _05830_ (
  .A1(_00887_),
  .A2(_00888_),
  .ZN(_00889_)
);

NAND2_X1 _05831_ (
  .A1(_00889_),
  .A2(_00857_),
  .ZN(_00890_)
);

NAND2_X1 _05832_ (
  .A1(_00870_),
  .A2(\sresult[2][2] ),
  .ZN(_00891_)
);

NAND2_X1 _05833_ (
  .A1(_00890_),
  .A2(_00891_),
  .ZN(_00026_)
);

NAND2_X1 _05834_ (
  .A1(_00865_),
  .A2(\sresult[1][3] ),
  .ZN(_00892_)
);

NAND2_X1 _05835_ (
  .A1(_00854_),
  .A2(din_67[3]),
  .ZN(_00893_)
);

NAND2_X1 _05836_ (
  .A1(_00892_),
  .A2(_00893_),
  .ZN(_00894_)
);

NAND2_X1 _05837_ (
  .A1(_00894_),
  .A2(_00857_),
  .ZN(_00895_)
);

NAND2_X1 _05838_ (
  .A1(_00870_),
  .A2(\sresult[2][3] ),
  .ZN(_00896_)
);

NAND2_X1 _05839_ (
  .A1(_00895_),
  .A2(_00896_),
  .ZN(_00027_)
);

NAND2_X1 _05840_ (
  .A1(_00865_),
  .A2(\sresult[1][4] ),
  .ZN(_00897_)
);

NAND2_X1 _05841_ (
  .A1(_00854_),
  .A2(din_67[4]),
  .ZN(_00898_)
);

NAND2_X1 _05842_ (
  .A1(_00897_),
  .A2(_00898_),
  .ZN(_00899_)
);

NAND2_X1 _05843_ (
  .A1(_00899_),
  .A2(_00857_),
  .ZN(_00900_)
);

NAND2_X1 _05844_ (
  .A1(_00870_),
  .A2(\sresult[2][4] ),
  .ZN(_00901_)
);

NAND2_X1 _05845_ (
  .A1(_00900_),
  .A2(_00901_),
  .ZN(_00028_)
);

NAND2_X1 _05846_ (
  .A1(_00865_),
  .A2(\sresult[1][5] ),
  .ZN(_00902_)
);

NAND2_X1 _05847_ (
  .A1(_00854_),
  .A2(din_67[5]),
  .ZN(_00903_)
);

NAND2_X1 _05848_ (
  .A1(_00902_),
  .A2(_00903_),
  .ZN(_00904_)
);

NAND2_X1 _05849_ (
  .A1(_00904_),
  .A2(_00857_),
  .ZN(_00905_)
);

NAND2_X1 _05850_ (
  .A1(_00870_),
  .A2(\sresult[2][5] ),
  .ZN(_00906_)
);

NAND2_X1 _05851_ (
  .A1(_00905_),
  .A2(_00906_),
  .ZN(_00029_)
);

NAND2_X1 _05852_ (
  .A1(_00865_),
  .A2(\sresult[1][6] ),
  .ZN(_00907_)
);

BUF_X4 _05853_ (
  .A(_00803_),
  .Z(_00908_)
);

NAND2_X1 _05854_ (
  .A1(_00908_),
  .A2(din_67[6]),
  .ZN(_00909_)
);

NAND2_X1 _05855_ (
  .A1(_00907_),
  .A2(_00909_),
  .ZN(_00910_)
);

BUF_X8 _05856_ (
  .A(_00771_),
  .Z(_00911_)
);

BUF_X4 _05857_ (
  .A(_00911_),
  .Z(_00912_)
);

BUF_X2 _05858_ (
  .A(_00912_),
  .Z(_00913_)
);

NAND2_X1 _05859_ (
  .A1(_00910_),
  .A2(_00913_),
  .ZN(_00914_)
);

NAND2_X1 _05860_ (
  .A1(_00870_),
  .A2(\sresult[2][6] ),
  .ZN(_00915_)
);

NAND2_X1 _05861_ (
  .A1(_00914_),
  .A2(_00915_),
  .ZN(_00030_)
);

NAND2_X1 _05862_ (
  .A1(_00865_),
  .A2(\sresult[1][7] ),
  .ZN(_00916_)
);

NAND2_X1 _05863_ (
  .A1(_00908_),
  .A2(din_67[7]),
  .ZN(_00917_)
);

NAND2_X1 _05864_ (
  .A1(_00916_),
  .A2(_00917_),
  .ZN(_00918_)
);

NAND2_X1 _05865_ (
  .A1(_00918_),
  .A2(_00913_),
  .ZN(_00919_)
);

NAND2_X1 _05866_ (
  .A1(_00870_),
  .A2(\sresult[2][7] ),
  .ZN(_00920_)
);

NAND2_X1 _05867_ (
  .A1(_00919_),
  .A2(_00920_),
  .ZN(_00031_)
);

BUF_X4 _05868_ (
  .A(_00814_),
  .Z(_00921_)
);

NAND2_X1 _05869_ (
  .A1(_00921_),
  .A2(\sresult[1][8] ),
  .ZN(_00922_)
);

NAND2_X1 _05870_ (
  .A1(_00908_),
  .A2(din_67[8]),
  .ZN(_00923_)
);

NAND2_X1 _05871_ (
  .A1(_00922_),
  .A2(_00923_),
  .ZN(_00924_)
);

NAND2_X1 _05872_ (
  .A1(_00924_),
  .A2(_00913_),
  .ZN(_00925_)
);

CLKBUF_X2 _05873_ (
  .A(_00820_),
  .Z(_00926_)
);

NAND2_X1 _05874_ (
  .A1(_00926_),
  .A2(\sresult[2][8] ),
  .ZN(_00927_)
);

NAND2_X1 _05875_ (
  .A1(_00925_),
  .A2(_00927_),
  .ZN(_00032_)
);

NAND2_X1 _05876_ (
  .A1(_00921_),
  .A2(\sresult[1][9] ),
  .ZN(_00928_)
);

NAND2_X1 _05877_ (
  .A1(_00908_),
  .A2(din_67[9]),
  .ZN(_00929_)
);

NAND2_X1 _05878_ (
  .A1(_00928_),
  .A2(_00929_),
  .ZN(_00930_)
);

NAND2_X1 _05879_ (
  .A1(_00930_),
  .A2(_00913_),
  .ZN(_00931_)
);

NAND2_X1 _05880_ (
  .A1(_00926_),
  .A2(\sresult[2][9] ),
  .ZN(_00932_)
);

NAND2_X1 _05881_ (
  .A1(_00931_),
  .A2(_00932_),
  .ZN(_00033_)
);

NAND2_X1 _05882_ (
  .A1(_00921_),
  .A2(\sresult[1][10] ),
  .ZN(_00933_)
);

NAND2_X1 _05883_ (
  .A1(_00908_),
  .A2(din_67[10]),
  .ZN(_00934_)
);

NAND2_X1 _05884_ (
  .A1(_00933_),
  .A2(_00934_),
  .ZN(_00935_)
);

NAND2_X1 _05885_ (
  .A1(_00935_),
  .A2(_00913_),
  .ZN(_00936_)
);

NAND2_X1 _05886_ (
  .A1(_00926_),
  .A2(\sresult[2][10] ),
  .ZN(_00937_)
);

NAND2_X1 _05887_ (
  .A1(_00936_),
  .A2(_00937_),
  .ZN(_00034_)
);

NAND2_X1 _05888_ (
  .A1(_00921_),
  .A2(\sresult[1][11] ),
  .ZN(_00938_)
);

NAND2_X1 _05889_ (
  .A1(_00908_),
  .A2(din_67[11]),
  .ZN(_00939_)
);

NAND2_X1 _05890_ (
  .A1(_00938_),
  .A2(_00939_),
  .ZN(_00940_)
);

NAND2_X1 _05891_ (
  .A1(_00940_),
  .A2(_00913_),
  .ZN(_00941_)
);

NAND2_X1 _05892_ (
  .A1(_00926_),
  .A2(\sresult[2][11] ),
  .ZN(_00942_)
);

NAND2_X1 _05893_ (
  .A1(_00941_),
  .A2(_00942_),
  .ZN(_00035_)
);

NAND2_X1 _05894_ (
  .A1(_00921_),
  .A2(\sresult[2][0] ),
  .ZN(_00943_)
);

NAND2_X1 _05895_ (
  .A1(_00908_),
  .A2(din_57[0]),
  .ZN(_00944_)
);

NAND2_X1 _05896_ (
  .A1(_00943_),
  .A2(_00944_),
  .ZN(_00945_)
);

NAND2_X1 _05897_ (
  .A1(_00945_),
  .A2(_00913_),
  .ZN(_00946_)
);

NAND2_X1 _05898_ (
  .A1(_00926_),
  .A2(\sresult[3][0] ),
  .ZN(_00947_)
);

NAND2_X1 _05899_ (
  .A1(_00946_),
  .A2(_00947_),
  .ZN(_00036_)
);

NAND2_X1 _05900_ (
  .A1(_00921_),
  .A2(\sresult[2][1] ),
  .ZN(_00948_)
);

NAND2_X1 _05901_ (
  .A1(_00908_),
  .A2(din_57[1]),
  .ZN(_00949_)
);

NAND2_X1 _05902_ (
  .A1(_00948_),
  .A2(_00949_),
  .ZN(_00950_)
);

NAND2_X1 _05903_ (
  .A1(_00950_),
  .A2(_00913_),
  .ZN(_00951_)
);

NAND2_X1 _05904_ (
  .A1(_00926_),
  .A2(\sresult[3][1] ),
  .ZN(_00952_)
);

NAND2_X1 _05905_ (
  .A1(_00951_),
  .A2(_00952_),
  .ZN(_00037_)
);

NAND2_X1 _05906_ (
  .A1(_00921_),
  .A2(\sresult[2][2] ),
  .ZN(_00953_)
);

NAND2_X1 _05907_ (
  .A1(_00908_),
  .A2(din_57[2]),
  .ZN(_00954_)
);

NAND2_X1 _05908_ (
  .A1(_00953_),
  .A2(_00954_),
  .ZN(_00955_)
);

NAND2_X1 _05909_ (
  .A1(_00955_),
  .A2(_00913_),
  .ZN(_00956_)
);

NAND2_X1 _05910_ (
  .A1(_00926_),
  .A2(\sresult[3][2] ),
  .ZN(_00957_)
);

NAND2_X1 _05911_ (
  .A1(_00956_),
  .A2(_00957_),
  .ZN(_00038_)
);

NAND2_X1 _05912_ (
  .A1(_00921_),
  .A2(\sresult[2][3] ),
  .ZN(_00958_)
);

NAND2_X1 _05913_ (
  .A1(_00908_),
  .A2(din_57[3]),
  .ZN(_00959_)
);

NAND2_X1 _05914_ (
  .A1(_00958_),
  .A2(_00959_),
  .ZN(_00960_)
);

NAND2_X1 _05915_ (
  .A1(_00960_),
  .A2(_00913_),
  .ZN(_00961_)
);

NAND2_X1 _05916_ (
  .A1(_00926_),
  .A2(\sresult[3][3] ),
  .ZN(_00962_)
);

NAND2_X1 _05917_ (
  .A1(_00961_),
  .A2(_00962_),
  .ZN(_00039_)
);

NAND2_X1 _05918_ (
  .A1(_00921_),
  .A2(\sresult[2][4] ),
  .ZN(_00963_)
);

BUF_X4 _05919_ (
  .A(_00803_),
  .Z(_00964_)
);

NAND2_X1 _05920_ (
  .A1(_00964_),
  .A2(din_57[4]),
  .ZN(_00965_)
);

NAND2_X1 _05921_ (
  .A1(_00963_),
  .A2(_00965_),
  .ZN(_00966_)
);

BUF_X2 _05922_ (
  .A(_00912_),
  .Z(_00967_)
);

NAND2_X1 _05923_ (
  .A1(_00966_),
  .A2(_00967_),
  .ZN(_00968_)
);

NAND2_X1 _05924_ (
  .A1(_00926_),
  .A2(\sresult[3][4] ),
  .ZN(_00969_)
);

NAND2_X1 _05925_ (
  .A1(_00968_),
  .A2(_00969_),
  .ZN(_00040_)
);

NAND2_X1 _05926_ (
  .A1(_00921_),
  .A2(\sresult[2][5] ),
  .ZN(_00970_)
);

NAND2_X1 _05927_ (
  .A1(_00964_),
  .A2(din_57[5]),
  .ZN(_00971_)
);

NAND2_X1 _05928_ (
  .A1(_00970_),
  .A2(_00971_),
  .ZN(_00972_)
);

NAND2_X1 _05929_ (
  .A1(_00972_),
  .A2(_00967_),
  .ZN(_00973_)
);

NAND2_X1 _05930_ (
  .A1(_00926_),
  .A2(\sresult[3][5] ),
  .ZN(_00974_)
);

NAND2_X1 _05931_ (
  .A1(_00973_),
  .A2(_00974_),
  .ZN(_00041_)
);

BUF_X8 _05932_ (
  .A(_00799_),
  .Z(_00975_)
);

BUF_X4 _05933_ (
  .A(_00975_),
  .Z(_00976_)
);

NAND2_X1 _05934_ (
  .A1(_00976_),
  .A2(\sresult[2][6] ),
  .ZN(_00977_)
);

NAND2_X1 _05935_ (
  .A1(_00964_),
  .A2(din_57[6]),
  .ZN(_00978_)
);

NAND2_X1 _05936_ (
  .A1(_00977_),
  .A2(_00978_),
  .ZN(_00979_)
);

NAND2_X1 _05937_ (
  .A1(_00979_),
  .A2(_00967_),
  .ZN(_00980_)
);

CLKBUF_X2 _05938_ (
  .A(_00820_),
  .Z(_00981_)
);

NAND2_X1 _05939_ (
  .A1(_00981_),
  .A2(\sresult[3][6] ),
  .ZN(_00982_)
);

NAND2_X1 _05940_ (
  .A1(_00980_),
  .A2(_00982_),
  .ZN(_00042_)
);

NAND2_X1 _05941_ (
  .A1(_00976_),
  .A2(\sresult[2][7] ),
  .ZN(_00983_)
);

NAND2_X1 _05942_ (
  .A1(_00964_),
  .A2(din_57[7]),
  .ZN(_00984_)
);

NAND2_X1 _05943_ (
  .A1(_00983_),
  .A2(_00984_),
  .ZN(_00985_)
);

NAND2_X1 _05944_ (
  .A1(_00985_),
  .A2(_00967_),
  .ZN(_00986_)
);

NAND2_X1 _05945_ (
  .A1(_00981_),
  .A2(\sresult[3][7] ),
  .ZN(_00987_)
);

NAND2_X1 _05946_ (
  .A1(_00986_),
  .A2(_00987_),
  .ZN(_00043_)
);

NAND2_X1 _05947_ (
  .A1(_00976_),
  .A2(\sresult[2][8] ),
  .ZN(_00988_)
);

NAND2_X1 _05948_ (
  .A1(_00964_),
  .A2(din_57[8]),
  .ZN(_00989_)
);

NAND2_X1 _05949_ (
  .A1(_00988_),
  .A2(_00989_),
  .ZN(_00990_)
);

NAND2_X1 _05950_ (
  .A1(_00990_),
  .A2(_00967_),
  .ZN(_00991_)
);

NAND2_X1 _05951_ (
  .A1(_00981_),
  .A2(\sresult[3][8] ),
  .ZN(_00992_)
);

NAND2_X1 _05952_ (
  .A1(_00991_),
  .A2(_00992_),
  .ZN(_00044_)
);

NAND2_X1 _05953_ (
  .A1(_00976_),
  .A2(\sresult[2][9] ),
  .ZN(_00993_)
);

NAND2_X1 _05954_ (
  .A1(_00964_),
  .A2(din_57[9]),
  .ZN(_00994_)
);

NAND2_X1 _05955_ (
  .A1(_00993_),
  .A2(_00994_),
  .ZN(_00995_)
);

NAND2_X1 _05956_ (
  .A1(_00995_),
  .A2(_00967_),
  .ZN(_00996_)
);

NAND2_X1 _05957_ (
  .A1(_00981_),
  .A2(\sresult[3][9] ),
  .ZN(_00997_)
);

NAND2_X1 _05958_ (
  .A1(_00996_),
  .A2(_00997_),
  .ZN(_00045_)
);

NAND2_X1 _05959_ (
  .A1(_00976_),
  .A2(\sresult[2][10] ),
  .ZN(_00998_)
);

NAND2_X1 _05960_ (
  .A1(_00964_),
  .A2(din_57[10]),
  .ZN(_00999_)
);

NAND2_X1 _05961_ (
  .A1(_00998_),
  .A2(_00999_),
  .ZN(_01000_)
);

NAND2_X1 _05962_ (
  .A1(_01000_),
  .A2(_00967_),
  .ZN(_01001_)
);

NAND2_X1 _05963_ (
  .A1(_00981_),
  .A2(\sresult[3][10] ),
  .ZN(_01002_)
);

NAND2_X1 _05964_ (
  .A1(_01001_),
  .A2(_01002_),
  .ZN(_00046_)
);

NAND2_X1 _05965_ (
  .A1(_00976_),
  .A2(\sresult[2][11] ),
  .ZN(_01003_)
);

NAND2_X1 _05966_ (
  .A1(_00964_),
  .A2(din_57[11]),
  .ZN(_01004_)
);

NAND2_X1 _05967_ (
  .A1(_01003_),
  .A2(_01004_),
  .ZN(_01005_)
);

NAND2_X1 _05968_ (
  .A1(_01005_),
  .A2(_00967_),
  .ZN(_01006_)
);

NAND2_X1 _05969_ (
  .A1(_00981_),
  .A2(\sresult[3][11] ),
  .ZN(_01007_)
);

NAND2_X1 _05970_ (
  .A1(_01006_),
  .A2(_01007_),
  .ZN(_00047_)
);

NAND2_X1 _05971_ (
  .A1(_00976_),
  .A2(\sresult[3][0] ),
  .ZN(_01008_)
);

NAND2_X1 _05972_ (
  .A1(_00964_),
  .A2(din_66[0]),
  .ZN(_01009_)
);

NAND2_X1 _05973_ (
  .A1(_01008_),
  .A2(_01009_),
  .ZN(_01010_)
);

NAND2_X1 _05974_ (
  .A1(_01010_),
  .A2(_00967_),
  .ZN(_01011_)
);

NAND2_X1 _05975_ (
  .A1(_00981_),
  .A2(\sresult[4][0] ),
  .ZN(_01012_)
);

NAND2_X1 _05976_ (
  .A1(_01011_),
  .A2(_01012_),
  .ZN(_00048_)
);

NAND2_X1 _05977_ (
  .A1(_00976_),
  .A2(\sresult[3][1] ),
  .ZN(_01013_)
);

NAND2_X1 _05978_ (
  .A1(_00964_),
  .A2(din_66[1]),
  .ZN(_01014_)
);

NAND2_X1 _05979_ (
  .A1(_01013_),
  .A2(_01014_),
  .ZN(_01015_)
);

NAND2_X1 _05980_ (
  .A1(_01015_),
  .A2(_00967_),
  .ZN(_01016_)
);

NAND2_X1 _05981_ (
  .A1(_00981_),
  .A2(\sresult[4][1] ),
  .ZN(_01017_)
);

NAND2_X1 _05982_ (
  .A1(_01016_),
  .A2(_01017_),
  .ZN(_00049_)
);

NAND2_X1 _05983_ (
  .A1(_00976_),
  .A2(\sresult[3][2] ),
  .ZN(_01018_)
);

BUF_X8 _05984_ (
  .A(_00770_),
  .Z(_01019_)
);

BUF_X4 _05985_ (
  .A(_01019_),
  .Z(_01020_)
);

NAND2_X1 _05986_ (
  .A1(_01020_),
  .A2(din_66[2]),
  .ZN(_01021_)
);

NAND2_X1 _05987_ (
  .A1(_01018_),
  .A2(_01021_),
  .ZN(_01022_)
);

BUF_X2 _05988_ (
  .A(_00912_),
  .Z(_01023_)
);

NAND2_X1 _05989_ (
  .A1(_01022_),
  .A2(_01023_),
  .ZN(_01024_)
);

NAND2_X1 _05990_ (
  .A1(_00981_),
  .A2(\sresult[4][2] ),
  .ZN(_01025_)
);

NAND2_X1 _05991_ (
  .A1(_01024_),
  .A2(_01025_),
  .ZN(_00050_)
);

NAND2_X1 _05992_ (
  .A1(_00976_),
  .A2(\sresult[3][3] ),
  .ZN(_01026_)
);

NAND2_X1 _05993_ (
  .A1(_01020_),
  .A2(din_66[3]),
  .ZN(_01027_)
);

NAND2_X1 _05994_ (
  .A1(_01026_),
  .A2(_01027_),
  .ZN(_01028_)
);

NAND2_X1 _05995_ (
  .A1(_01028_),
  .A2(_01023_),
  .ZN(_01029_)
);

NAND2_X1 _05996_ (
  .A1(_00981_),
  .A2(\sresult[4][3] ),
  .ZN(_01030_)
);

NAND2_X1 _05997_ (
  .A1(_01029_),
  .A2(_01030_),
  .ZN(_00051_)
);

BUF_X4 _05998_ (
  .A(_00975_),
  .Z(_01031_)
);

NAND2_X1 _05999_ (
  .A1(_01031_),
  .A2(\sresult[3][4] ),
  .ZN(_01032_)
);

NAND2_X1 _06000_ (
  .A1(_01020_),
  .A2(din_66[4]),
  .ZN(_01033_)
);

NAND2_X1 _06001_ (
  .A1(_01032_),
  .A2(_01033_),
  .ZN(_01034_)
);

NAND2_X1 _06002_ (
  .A1(_01034_),
  .A2(_01023_),
  .ZN(_01035_)
);

BUF_X4 _06003_ (
  .A(_00810_),
  .Z(_01036_)
);

CLKBUF_X2 _06004_ (
  .A(_01036_),
  .Z(_01037_)
);

NAND2_X1 _06005_ (
  .A1(_01037_),
  .A2(\sresult[4][4] ),
  .ZN(_01038_)
);

NAND2_X1 _06006_ (
  .A1(_01035_),
  .A2(_01038_),
  .ZN(_00052_)
);

NAND2_X1 _06007_ (
  .A1(_01031_),
  .A2(\sresult[3][5] ),
  .ZN(_01039_)
);

NAND2_X1 _06008_ (
  .A1(_01020_),
  .A2(din_66[5]),
  .ZN(_01040_)
);

NAND2_X1 _06009_ (
  .A1(_01039_),
  .A2(_01040_),
  .ZN(_01041_)
);

NAND2_X1 _06010_ (
  .A1(_01041_),
  .A2(_01023_),
  .ZN(_01042_)
);

NAND2_X1 _06011_ (
  .A1(_01037_),
  .A2(\sresult[4][5] ),
  .ZN(_01043_)
);

NAND2_X1 _06012_ (
  .A1(_01042_),
  .A2(_01043_),
  .ZN(_00053_)
);

NAND2_X1 _06013_ (
  .A1(_01031_),
  .A2(\sresult[3][6] ),
  .ZN(_01044_)
);

NAND2_X1 _06014_ (
  .A1(_01020_),
  .A2(din_66[6]),
  .ZN(_01045_)
);

NAND2_X1 _06015_ (
  .A1(_01044_),
  .A2(_01045_),
  .ZN(_01046_)
);

NAND2_X1 _06016_ (
  .A1(_01046_),
  .A2(_01023_),
  .ZN(_01047_)
);

NAND2_X1 _06017_ (
  .A1(_01037_),
  .A2(\sresult[4][6] ),
  .ZN(_01048_)
);

NAND2_X1 _06018_ (
  .A1(_01047_),
  .A2(_01048_),
  .ZN(_00054_)
);

NAND2_X1 _06019_ (
  .A1(_01031_),
  .A2(\sresult[3][7] ),
  .ZN(_01049_)
);

NAND2_X1 _06020_ (
  .A1(_01020_),
  .A2(din_66[7]),
  .ZN(_01050_)
);

NAND2_X1 _06021_ (
  .A1(_01049_),
  .A2(_01050_),
  .ZN(_01051_)
);

NAND2_X1 _06022_ (
  .A1(_01051_),
  .A2(_01023_),
  .ZN(_01052_)
);

NAND2_X1 _06023_ (
  .A1(_01037_),
  .A2(\sresult[4][7] ),
  .ZN(_01053_)
);

NAND2_X1 _06024_ (
  .A1(_01052_),
  .A2(_01053_),
  .ZN(_00055_)
);

NAND2_X1 _06025_ (
  .A1(_01031_),
  .A2(\sresult[3][8] ),
  .ZN(_01054_)
);

NAND2_X1 _06026_ (
  .A1(_01020_),
  .A2(din_66[8]),
  .ZN(_01055_)
);

NAND2_X1 _06027_ (
  .A1(_01054_),
  .A2(_01055_),
  .ZN(_01056_)
);

NAND2_X1 _06028_ (
  .A1(_01056_),
  .A2(_01023_),
  .ZN(_01057_)
);

NAND2_X1 _06029_ (
  .A1(_01037_),
  .A2(\sresult[4][8] ),
  .ZN(_01058_)
);

NAND2_X1 _06030_ (
  .A1(_01057_),
  .A2(_01058_),
  .ZN(_00056_)
);

NAND2_X1 _06031_ (
  .A1(_01031_),
  .A2(\sresult[3][9] ),
  .ZN(_01059_)
);

NAND2_X1 _06032_ (
  .A1(_01020_),
  .A2(din_66[9]),
  .ZN(_01060_)
);

NAND2_X1 _06033_ (
  .A1(_01059_),
  .A2(_01060_),
  .ZN(_01061_)
);

NAND2_X1 _06034_ (
  .A1(_01061_),
  .A2(_01023_),
  .ZN(_01062_)
);

NAND2_X1 _06035_ (
  .A1(_01037_),
  .A2(\sresult[4][9] ),
  .ZN(_01063_)
);

NAND2_X1 _06036_ (
  .A1(_01062_),
  .A2(_01063_),
  .ZN(_00057_)
);

NAND2_X1 _06037_ (
  .A1(_01031_),
  .A2(\sresult[3][10] ),
  .ZN(_01064_)
);

NAND2_X1 _06038_ (
  .A1(_01020_),
  .A2(din_66[10]),
  .ZN(_01065_)
);

NAND2_X1 _06039_ (
  .A1(_01064_),
  .A2(_01065_),
  .ZN(_01066_)
);

NAND2_X1 _06040_ (
  .A1(_01066_),
  .A2(_01023_),
  .ZN(_01067_)
);

NAND2_X1 _06041_ (
  .A1(_01037_),
  .A2(\sresult[4][10] ),
  .ZN(_01068_)
);

NAND2_X1 _06042_ (
  .A1(_01067_),
  .A2(_01068_),
  .ZN(_00058_)
);

NAND2_X1 _06043_ (
  .A1(_01031_),
  .A2(\sresult[3][11] ),
  .ZN(_01069_)
);

NAND2_X1 _06044_ (
  .A1(_01020_),
  .A2(din_66[11]),
  .ZN(_01070_)
);

NAND2_X1 _06045_ (
  .A1(_01069_),
  .A2(_01070_),
  .ZN(_01071_)
);

NAND2_X1 _06046_ (
  .A1(_01071_),
  .A2(_01023_),
  .ZN(_01072_)
);

NAND2_X1 _06047_ (
  .A1(_01037_),
  .A2(\sresult[4][11] ),
  .ZN(_01073_)
);

NAND2_X1 _06048_ (
  .A1(_01072_),
  .A2(_01073_),
  .ZN(_00059_)
);

NAND2_X1 _06049_ (
  .A1(_01031_),
  .A2(\sresult[4][0] ),
  .ZN(_01074_)
);

BUF_X4 _06050_ (
  .A(_01019_),
  .Z(_01075_)
);

NAND2_X1 _06051_ (
  .A1(_01075_),
  .A2(din_75[0]),
  .ZN(_01076_)
);

NAND2_X1 _06052_ (
  .A1(_01074_),
  .A2(_01076_),
  .ZN(_01077_)
);

BUF_X2 _06053_ (
  .A(_00912_),
  .Z(_01078_)
);

NAND2_X1 _06054_ (
  .A1(_01077_),
  .A2(_01078_),
  .ZN(_01079_)
);

NAND2_X1 _06055_ (
  .A1(_01037_),
  .A2(\sresult[5][0] ),
  .ZN(_01080_)
);

NAND2_X1 _06056_ (
  .A1(_01079_),
  .A2(_01080_),
  .ZN(_00060_)
);

NAND2_X1 _06057_ (
  .A1(_01031_),
  .A2(\sresult[4][1] ),
  .ZN(_01081_)
);

NAND2_X1 _06058_ (
  .A1(_01075_),
  .A2(din_75[1]),
  .ZN(_01082_)
);

NAND2_X1 _06059_ (
  .A1(_01081_),
  .A2(_01082_),
  .ZN(_01083_)
);

NAND2_X1 _06060_ (
  .A1(_01083_),
  .A2(_01078_),
  .ZN(_01084_)
);

NAND2_X1 _06061_ (
  .A1(_01037_),
  .A2(\sresult[5][1] ),
  .ZN(_01085_)
);

NAND2_X1 _06062_ (
  .A1(_01084_),
  .A2(_01085_),
  .ZN(_00061_)
);

BUF_X4 _06063_ (
  .A(_00975_),
  .Z(_01086_)
);

NAND2_X1 _06064_ (
  .A1(_01086_),
  .A2(\sresult[4][2] ),
  .ZN(_01087_)
);

NAND2_X1 _06065_ (
  .A1(_01075_),
  .A2(din_75[2]),
  .ZN(_01088_)
);

NAND2_X1 _06066_ (
  .A1(_01087_),
  .A2(_01088_),
  .ZN(_01089_)
);

NAND2_X1 _06067_ (
  .A1(_01089_),
  .A2(_01078_),
  .ZN(_01090_)
);

CLKBUF_X2 _06068_ (
  .A(_01036_),
  .Z(_01091_)
);

NAND2_X1 _06069_ (
  .A1(_01091_),
  .A2(\sresult[5][2] ),
  .ZN(_01092_)
);

NAND2_X1 _06070_ (
  .A1(_01090_),
  .A2(_01092_),
  .ZN(_00062_)
);

NAND2_X1 _06071_ (
  .A1(_01086_),
  .A2(\sresult[4][3] ),
  .ZN(_01093_)
);

NAND2_X1 _06072_ (
  .A1(_01075_),
  .A2(din_75[3]),
  .ZN(_01094_)
);

NAND2_X1 _06073_ (
  .A1(_01093_),
  .A2(_01094_),
  .ZN(_01095_)
);

NAND2_X1 _06074_ (
  .A1(_01095_),
  .A2(_01078_),
  .ZN(_01096_)
);

NAND2_X1 _06075_ (
  .A1(_01091_),
  .A2(\sresult[5][3] ),
  .ZN(_01097_)
);

NAND2_X1 _06076_ (
  .A1(_01096_),
  .A2(_01097_),
  .ZN(_00063_)
);

NAND2_X1 _06077_ (
  .A1(_01086_),
  .A2(\sresult[4][4] ),
  .ZN(_01098_)
);

NAND2_X1 _06078_ (
  .A1(_01075_),
  .A2(din_75[4]),
  .ZN(_01099_)
);

NAND2_X1 _06079_ (
  .A1(_01098_),
  .A2(_01099_),
  .ZN(_01100_)
);

NAND2_X1 _06080_ (
  .A1(_01100_),
  .A2(_01078_),
  .ZN(_01101_)
);

NAND2_X1 _06081_ (
  .A1(_01091_),
  .A2(\sresult[5][4] ),
  .ZN(_01102_)
);

NAND2_X1 _06082_ (
  .A1(_01101_),
  .A2(_01102_),
  .ZN(_00064_)
);

NAND2_X1 _06083_ (
  .A1(_01086_),
  .A2(\sresult[4][5] ),
  .ZN(_01103_)
);

NAND2_X1 _06084_ (
  .A1(_01075_),
  .A2(din_75[5]),
  .ZN(_01104_)
);

NAND2_X1 _06085_ (
  .A1(_01103_),
  .A2(_01104_),
  .ZN(_01105_)
);

NAND2_X1 _06086_ (
  .A1(_01105_),
  .A2(_01078_),
  .ZN(_01106_)
);

NAND2_X1 _06087_ (
  .A1(_01091_),
  .A2(\sresult[5][5] ),
  .ZN(_01107_)
);

NAND2_X1 _06088_ (
  .A1(_01106_),
  .A2(_01107_),
  .ZN(_00065_)
);

NAND2_X1 _06089_ (
  .A1(_01086_),
  .A2(\sresult[4][6] ),
  .ZN(_01108_)
);

NAND2_X1 _06090_ (
  .A1(_01075_),
  .A2(din_75[6]),
  .ZN(_01109_)
);

NAND2_X1 _06091_ (
  .A1(_01108_),
  .A2(_01109_),
  .ZN(_01110_)
);

NAND2_X1 _06092_ (
  .A1(_01110_),
  .A2(_01078_),
  .ZN(_01111_)
);

NAND2_X1 _06093_ (
  .A1(_01091_),
  .A2(\sresult[5][6] ),
  .ZN(_01112_)
);

NAND2_X1 _06094_ (
  .A1(_01111_),
  .A2(_01112_),
  .ZN(_00066_)
);

NAND2_X1 _06095_ (
  .A1(_01086_),
  .A2(\sresult[4][7] ),
  .ZN(_01113_)
);

NAND2_X1 _06096_ (
  .A1(_01075_),
  .A2(din_75[7]),
  .ZN(_01114_)
);

NAND2_X1 _06097_ (
  .A1(_01113_),
  .A2(_01114_),
  .ZN(_01115_)
);

NAND2_X1 _06098_ (
  .A1(_01115_),
  .A2(_01078_),
  .ZN(_01116_)
);

NAND2_X1 _06099_ (
  .A1(_01091_),
  .A2(\sresult[5][7] ),
  .ZN(_01117_)
);

NAND2_X1 _06100_ (
  .A1(_01116_),
  .A2(_01117_),
  .ZN(_00067_)
);

NAND2_X1 _06101_ (
  .A1(_01086_),
  .A2(\sresult[4][8] ),
  .ZN(_01118_)
);

NAND2_X1 _06102_ (
  .A1(_01075_),
  .A2(din_75[8]),
  .ZN(_01119_)
);

NAND2_X1 _06103_ (
  .A1(_01118_),
  .A2(_01119_),
  .ZN(_01120_)
);

NAND2_X1 _06104_ (
  .A1(_01120_),
  .A2(_01078_),
  .ZN(_01121_)
);

NAND2_X1 _06105_ (
  .A1(_01091_),
  .A2(\sresult[5][8] ),
  .ZN(_01122_)
);

NAND2_X1 _06106_ (
  .A1(_01121_),
  .A2(_01122_),
  .ZN(_00068_)
);

NAND2_X1 _06107_ (
  .A1(_01086_),
  .A2(\sresult[4][9] ),
  .ZN(_01123_)
);

NAND2_X1 _06108_ (
  .A1(_01075_),
  .A2(din_75[9]),
  .ZN(_01124_)
);

NAND2_X1 _06109_ (
  .A1(_01123_),
  .A2(_01124_),
  .ZN(_01125_)
);

NAND2_X1 _06110_ (
  .A1(_01125_),
  .A2(_01078_),
  .ZN(_01126_)
);

NAND2_X1 _06111_ (
  .A1(_01091_),
  .A2(\sresult[5][9] ),
  .ZN(_01127_)
);

NAND2_X1 _06112_ (
  .A1(_01126_),
  .A2(_01127_),
  .ZN(_00069_)
);

NAND2_X1 _06113_ (
  .A1(_01086_),
  .A2(\sresult[4][10] ),
  .ZN(_01128_)
);

BUF_X4 _06114_ (
  .A(_01019_),
  .Z(_01129_)
);

NAND2_X1 _06115_ (
  .A1(_01129_),
  .A2(din_75[10]),
  .ZN(_01130_)
);

NAND2_X1 _06116_ (
  .A1(_01128_),
  .A2(_01130_),
  .ZN(_01131_)
);

BUF_X2 _06117_ (
  .A(_00912_),
  .Z(_01132_)
);

NAND2_X1 _06118_ (
  .A1(_01131_),
  .A2(_01132_),
  .ZN(_01133_)
);

NAND2_X1 _06119_ (
  .A1(_01091_),
  .A2(\sresult[5][10] ),
  .ZN(_01134_)
);

NAND2_X1 _06120_ (
  .A1(_01133_),
  .A2(_01134_),
  .ZN(_00070_)
);

NAND2_X1 _06121_ (
  .A1(_01086_),
  .A2(\sresult[4][11] ),
  .ZN(_01135_)
);

NAND2_X1 _06122_ (
  .A1(_01129_),
  .A2(din_75[11]),
  .ZN(_01136_)
);

NAND2_X1 _06123_ (
  .A1(_01135_),
  .A2(_01136_),
  .ZN(_01137_)
);

NAND2_X1 _06124_ (
  .A1(_01137_),
  .A2(_01132_),
  .ZN(_01138_)
);

NAND2_X1 _06125_ (
  .A1(_01091_),
  .A2(\sresult[5][11] ),
  .ZN(_01139_)
);

NAND2_X1 _06126_ (
  .A1(_01138_),
  .A2(_01139_),
  .ZN(_00071_)
);

BUF_X4 _06127_ (
  .A(_00975_),
  .Z(_01140_)
);

NAND2_X1 _06128_ (
  .A1(_01140_),
  .A2(\sresult[5][0] ),
  .ZN(_01141_)
);

NAND2_X1 _06129_ (
  .A1(_01129_),
  .A2(din_74[0]),
  .ZN(_01142_)
);

NAND2_X1 _06130_ (
  .A1(_01141_),
  .A2(_01142_),
  .ZN(_01143_)
);

NAND2_X1 _06131_ (
  .A1(_01143_),
  .A2(_01132_),
  .ZN(_01144_)
);

CLKBUF_X2 _06132_ (
  .A(_01036_),
  .Z(_01145_)
);

NAND2_X1 _06133_ (
  .A1(_01145_),
  .A2(\sresult[6][0] ),
  .ZN(_01146_)
);

NAND2_X1 _06134_ (
  .A1(_01144_),
  .A2(_01146_),
  .ZN(_00072_)
);

NAND2_X1 _06135_ (
  .A1(_01140_),
  .A2(\sresult[5][1] ),
  .ZN(_01147_)
);

NAND2_X1 _06136_ (
  .A1(_01129_),
  .A2(din_74[1]),
  .ZN(_01148_)
);

NAND2_X1 _06137_ (
  .A1(_01147_),
  .A2(_01148_),
  .ZN(_01149_)
);

NAND2_X1 _06138_ (
  .A1(_01149_),
  .A2(_01132_),
  .ZN(_01150_)
);

NAND2_X1 _06139_ (
  .A1(_01145_),
  .A2(\sresult[6][1] ),
  .ZN(_01151_)
);

NAND2_X1 _06140_ (
  .A1(_01150_),
  .A2(_01151_),
  .ZN(_00073_)
);

NAND2_X1 _06141_ (
  .A1(_01140_),
  .A2(\sresult[5][2] ),
  .ZN(_01152_)
);

NAND2_X1 _06142_ (
  .A1(_01129_),
  .A2(din_74[2]),
  .ZN(_01153_)
);

NAND2_X1 _06143_ (
  .A1(_01152_),
  .A2(_01153_),
  .ZN(_01154_)
);

NAND2_X1 _06144_ (
  .A1(_01154_),
  .A2(_01132_),
  .ZN(_01155_)
);

NAND2_X1 _06145_ (
  .A1(_01145_),
  .A2(\sresult[6][2] ),
  .ZN(_01156_)
);

NAND2_X1 _06146_ (
  .A1(_01155_),
  .A2(_01156_),
  .ZN(_00074_)
);

NAND2_X1 _06147_ (
  .A1(_01140_),
  .A2(\sresult[5][3] ),
  .ZN(_01157_)
);

NAND2_X1 _06148_ (
  .A1(_01129_),
  .A2(din_74[3]),
  .ZN(_01158_)
);

NAND2_X1 _06149_ (
  .A1(_01157_),
  .A2(_01158_),
  .ZN(_01159_)
);

NAND2_X1 _06150_ (
  .A1(_01159_),
  .A2(_01132_),
  .ZN(_01160_)
);

NAND2_X1 _06151_ (
  .A1(_01145_),
  .A2(\sresult[6][3] ),
  .ZN(_01161_)
);

NAND2_X1 _06152_ (
  .A1(_01160_),
  .A2(_01161_),
  .ZN(_00075_)
);

NAND2_X1 _06153_ (
  .A1(_01140_),
  .A2(\sresult[5][4] ),
  .ZN(_01162_)
);

NAND2_X1 _06154_ (
  .A1(_01129_),
  .A2(din_74[4]),
  .ZN(_01163_)
);

NAND2_X1 _06155_ (
  .A1(_01162_),
  .A2(_01163_),
  .ZN(_01164_)
);

NAND2_X1 _06156_ (
  .A1(_01164_),
  .A2(_01132_),
  .ZN(_01165_)
);

NAND2_X1 _06157_ (
  .A1(_01145_),
  .A2(\sresult[6][4] ),
  .ZN(_01166_)
);

NAND2_X1 _06158_ (
  .A1(_01165_),
  .A2(_01166_),
  .ZN(_00076_)
);

NAND2_X1 _06159_ (
  .A1(_01140_),
  .A2(\sresult[5][5] ),
  .ZN(_01167_)
);

NAND2_X1 _06160_ (
  .A1(_01129_),
  .A2(din_74[5]),
  .ZN(_01168_)
);

NAND2_X1 _06161_ (
  .A1(_01167_),
  .A2(_01168_),
  .ZN(_01169_)
);

NAND2_X1 _06162_ (
  .A1(_01169_),
  .A2(_01132_),
  .ZN(_01170_)
);

NAND2_X1 _06163_ (
  .A1(_01145_),
  .A2(\sresult[6][5] ),
  .ZN(_01171_)
);

NAND2_X1 _06164_ (
  .A1(_01170_),
  .A2(_01171_),
  .ZN(_00077_)
);

NAND2_X1 _06165_ (
  .A1(_01140_),
  .A2(\sresult[5][6] ),
  .ZN(_01172_)
);

NAND2_X1 _06166_ (
  .A1(_01129_),
  .A2(din_74[6]),
  .ZN(_01173_)
);

NAND2_X1 _06167_ (
  .A1(_01172_),
  .A2(_01173_),
  .ZN(_01174_)
);

NAND2_X1 _06168_ (
  .A1(_01174_),
  .A2(_01132_),
  .ZN(_01175_)
);

NAND2_X1 _06169_ (
  .A1(_01145_),
  .A2(\sresult[6][6] ),
  .ZN(_01176_)
);

NAND2_X1 _06170_ (
  .A1(_01175_),
  .A2(_01176_),
  .ZN(_00078_)
);

NAND2_X1 _06171_ (
  .A1(_01140_),
  .A2(\sresult[5][7] ),
  .ZN(_01177_)
);

NAND2_X1 _06172_ (
  .A1(_01129_),
  .A2(din_74[7]),
  .ZN(_01178_)
);

NAND2_X1 _06173_ (
  .A1(_01177_),
  .A2(_01178_),
  .ZN(_01179_)
);

NAND2_X1 _06174_ (
  .A1(_01179_),
  .A2(_01132_),
  .ZN(_01180_)
);

NAND2_X1 _06175_ (
  .A1(_01145_),
  .A2(\sresult[6][7] ),
  .ZN(_01181_)
);

NAND2_X1 _06176_ (
  .A1(_01180_),
  .A2(_01181_),
  .ZN(_00079_)
);

NAND2_X1 _06177_ (
  .A1(_01140_),
  .A2(\sresult[5][8] ),
  .ZN(_01182_)
);

BUF_X4 _06178_ (
  .A(_01019_),
  .Z(_01183_)
);

NAND2_X1 _06179_ (
  .A1(_01183_),
  .A2(din_74[8]),
  .ZN(_01184_)
);

NAND2_X1 _06180_ (
  .A1(_01182_),
  .A2(_01184_),
  .ZN(_01185_)
);

BUF_X2 _06181_ (
  .A(_00912_),
  .Z(_01186_)
);

NAND2_X1 _06182_ (
  .A1(_01185_),
  .A2(_01186_),
  .ZN(_01187_)
);

NAND2_X1 _06183_ (
  .A1(_01145_),
  .A2(\sresult[6][8] ),
  .ZN(_01188_)
);

NAND2_X1 _06184_ (
  .A1(_01187_),
  .A2(_01188_),
  .ZN(_00080_)
);

NAND2_X1 _06185_ (
  .A1(_01140_),
  .A2(\sresult[5][9] ),
  .ZN(_01189_)
);

NAND2_X1 _06186_ (
  .A1(_01183_),
  .A2(din_74[9]),
  .ZN(_01190_)
);

NAND2_X1 _06187_ (
  .A1(_01189_),
  .A2(_01190_),
  .ZN(_01191_)
);

NAND2_X1 _06188_ (
  .A1(_01191_),
  .A2(_01186_),
  .ZN(_01192_)
);

NAND2_X1 _06189_ (
  .A1(_01145_),
  .A2(\sresult[6][9] ),
  .ZN(_01193_)
);

NAND2_X1 _06190_ (
  .A1(_01192_),
  .A2(_01193_),
  .ZN(_00081_)
);

BUF_X4 _06191_ (
  .A(_00975_),
  .Z(_01194_)
);

NAND2_X1 _06192_ (
  .A1(_01194_),
  .A2(\sresult[5][10] ),
  .ZN(_01195_)
);

NAND2_X1 _06193_ (
  .A1(_01183_),
  .A2(din_74[10]),
  .ZN(_01196_)
);

NAND2_X1 _06194_ (
  .A1(_01195_),
  .A2(_01196_),
  .ZN(_01197_)
);

NAND2_X1 _06195_ (
  .A1(_01197_),
  .A2(_01186_),
  .ZN(_01198_)
);

CLKBUF_X2 _06196_ (
  .A(_01036_),
  .Z(_01199_)
);

NAND2_X1 _06197_ (
  .A1(_01199_),
  .A2(\sresult[6][10] ),
  .ZN(_01200_)
);

NAND2_X1 _06198_ (
  .A1(_01198_),
  .A2(_01200_),
  .ZN(_00082_)
);

NAND2_X1 _06199_ (
  .A1(_01194_),
  .A2(\sresult[5][11] ),
  .ZN(_01201_)
);

NAND2_X1 _06200_ (
  .A1(_01183_),
  .A2(din_74[11]),
  .ZN(_01202_)
);

NAND2_X1 _06201_ (
  .A1(_01201_),
  .A2(_01202_),
  .ZN(_01203_)
);

NAND2_X1 _06202_ (
  .A1(_01203_),
  .A2(_01186_),
  .ZN(_01204_)
);

NAND2_X1 _06203_ (
  .A1(_01199_),
  .A2(\sresult[6][11] ),
  .ZN(_01205_)
);

NAND2_X1 _06204_ (
  .A1(_01204_),
  .A2(_01205_),
  .ZN(_00083_)
);

NAND2_X1 _06205_ (
  .A1(_01194_),
  .A2(\sresult[6][0] ),
  .ZN(_01206_)
);

NAND2_X1 _06206_ (
  .A1(_01183_),
  .A2(din_65[0]),
  .ZN(_01207_)
);

NAND2_X1 _06207_ (
  .A1(_01206_),
  .A2(_01207_),
  .ZN(_01208_)
);

NAND2_X1 _06208_ (
  .A1(_01208_),
  .A2(_01186_),
  .ZN(_01209_)
);

NAND2_X1 _06209_ (
  .A1(_01199_),
  .A2(\sresult[7][0] ),
  .ZN(_01210_)
);

NAND2_X1 _06210_ (
  .A1(_01209_),
  .A2(_01210_),
  .ZN(_00084_)
);

NAND2_X1 _06211_ (
  .A1(_01194_),
  .A2(\sresult[6][1] ),
  .ZN(_01211_)
);

NAND2_X1 _06212_ (
  .A1(_01183_),
  .A2(din_65[1]),
  .ZN(_01212_)
);

NAND2_X1 _06213_ (
  .A1(_01211_),
  .A2(_01212_),
  .ZN(_01213_)
);

NAND2_X1 _06214_ (
  .A1(_01213_),
  .A2(_01186_),
  .ZN(_01214_)
);

NAND2_X1 _06215_ (
  .A1(_01199_),
  .A2(\sresult[7][1] ),
  .ZN(_01215_)
);

NAND2_X1 _06216_ (
  .A1(_01214_),
  .A2(_01215_),
  .ZN(_00085_)
);

NAND2_X1 _06217_ (
  .A1(_01194_),
  .A2(\sresult[6][2] ),
  .ZN(_01216_)
);

NAND2_X1 _06218_ (
  .A1(_01183_),
  .A2(din_65[2]),
  .ZN(_01217_)
);

NAND2_X1 _06219_ (
  .A1(_01216_),
  .A2(_01217_),
  .ZN(_01218_)
);

NAND2_X1 _06220_ (
  .A1(_01218_),
  .A2(_01186_),
  .ZN(_01219_)
);

NAND2_X1 _06221_ (
  .A1(_01199_),
  .A2(\sresult[7][2] ),
  .ZN(_01220_)
);

NAND2_X1 _06222_ (
  .A1(_01219_),
  .A2(_01220_),
  .ZN(_00086_)
);

NAND2_X1 _06223_ (
  .A1(_01194_),
  .A2(\sresult[6][3] ),
  .ZN(_01221_)
);

NAND2_X1 _06224_ (
  .A1(_01183_),
  .A2(din_65[3]),
  .ZN(_01222_)
);

NAND2_X1 _06225_ (
  .A1(_01221_),
  .A2(_01222_),
  .ZN(_01223_)
);

NAND2_X1 _06226_ (
  .A1(_01223_),
  .A2(_01186_),
  .ZN(_01224_)
);

NAND2_X1 _06227_ (
  .A1(_01199_),
  .A2(\sresult[7][3] ),
  .ZN(_01225_)
);

NAND2_X1 _06228_ (
  .A1(_01224_),
  .A2(_01225_),
  .ZN(_00087_)
);

NAND2_X1 _06229_ (
  .A1(_01194_),
  .A2(\sresult[6][4] ),
  .ZN(_01226_)
);

NAND2_X1 _06230_ (
  .A1(_01183_),
  .A2(din_65[4]),
  .ZN(_01227_)
);

NAND2_X1 _06231_ (
  .A1(_01226_),
  .A2(_01227_),
  .ZN(_01228_)
);

NAND2_X1 _06232_ (
  .A1(_01228_),
  .A2(_01186_),
  .ZN(_01229_)
);

NAND2_X1 _06233_ (
  .A1(_01199_),
  .A2(\sresult[7][4] ),
  .ZN(_01230_)
);

NAND2_X1 _06234_ (
  .A1(_01229_),
  .A2(_01230_),
  .ZN(_00088_)
);

NAND2_X1 _06235_ (
  .A1(_01194_),
  .A2(\sresult[6][5] ),
  .ZN(_01231_)
);

NAND2_X1 _06236_ (
  .A1(_01183_),
  .A2(din_65[5]),
  .ZN(_01232_)
);

NAND2_X1 _06237_ (
  .A1(_01231_),
  .A2(_01232_),
  .ZN(_01233_)
);

NAND2_X1 _06238_ (
  .A1(_01233_),
  .A2(_01186_),
  .ZN(_01234_)
);

NAND2_X1 _06239_ (
  .A1(_01199_),
  .A2(\sresult[7][5] ),
  .ZN(_01235_)
);

NAND2_X1 _06240_ (
  .A1(_01234_),
  .A2(_01235_),
  .ZN(_00089_)
);

NAND2_X1 _06241_ (
  .A1(_01194_),
  .A2(\sresult[6][6] ),
  .ZN(_01236_)
);

BUF_X4 _06242_ (
  .A(_01019_),
  .Z(_01237_)
);

NAND2_X1 _06243_ (
  .A1(_01237_),
  .A2(din_65[6]),
  .ZN(_01238_)
);

NAND2_X1 _06244_ (
  .A1(_01236_),
  .A2(_01238_),
  .ZN(_01239_)
);

BUF_X2 _06245_ (
  .A(_00912_),
  .Z(_01240_)
);

NAND2_X1 _06246_ (
  .A1(_01239_),
  .A2(_01240_),
  .ZN(_01241_)
);

NAND2_X1 _06247_ (
  .A1(_01199_),
  .A2(\sresult[7][6] ),
  .ZN(_01242_)
);

NAND2_X1 _06248_ (
  .A1(_01241_),
  .A2(_01242_),
  .ZN(_00090_)
);

NAND2_X1 _06249_ (
  .A1(_01194_),
  .A2(\sresult[6][7] ),
  .ZN(_01243_)
);

NAND2_X1 _06250_ (
  .A1(_01237_),
  .A2(din_65[7]),
  .ZN(_01244_)
);

NAND2_X1 _06251_ (
  .A1(_01243_),
  .A2(_01244_),
  .ZN(_01245_)
);

NAND2_X1 _06252_ (
  .A1(_01245_),
  .A2(_01240_),
  .ZN(_01246_)
);

NAND2_X1 _06253_ (
  .A1(_01199_),
  .A2(\sresult[7][7] ),
  .ZN(_01247_)
);

NAND2_X1 _06254_ (
  .A1(_01246_),
  .A2(_01247_),
  .ZN(_00091_)
);

BUF_X4 _06255_ (
  .A(_00975_),
  .Z(_01248_)
);

NAND2_X1 _06256_ (
  .A1(_01248_),
  .A2(\sresult[6][8] ),
  .ZN(_01249_)
);

NAND2_X1 _06257_ (
  .A1(_01237_),
  .A2(din_65[8]),
  .ZN(_01250_)
);

NAND2_X1 _06258_ (
  .A1(_01249_),
  .A2(_01250_),
  .ZN(_01251_)
);

NAND2_X1 _06259_ (
  .A1(_01251_),
  .A2(_01240_),
  .ZN(_01252_)
);

CLKBUF_X2 _06260_ (
  .A(_01036_),
  .Z(_01253_)
);

NAND2_X1 _06261_ (
  .A1(_01253_),
  .A2(\sresult[7][8] ),
  .ZN(_01254_)
);

NAND2_X1 _06262_ (
  .A1(_01252_),
  .A2(_01254_),
  .ZN(_00092_)
);

NAND2_X1 _06263_ (
  .A1(_01248_),
  .A2(\sresult[6][9] ),
  .ZN(_01255_)
);

NAND2_X1 _06264_ (
  .A1(_01237_),
  .A2(din_65[9]),
  .ZN(_01256_)
);

NAND2_X1 _06265_ (
  .A1(_01255_),
  .A2(_01256_),
  .ZN(_01257_)
);

NAND2_X1 _06266_ (
  .A1(_01257_),
  .A2(_01240_),
  .ZN(_01258_)
);

NAND2_X1 _06267_ (
  .A1(_01253_),
  .A2(\sresult[7][9] ),
  .ZN(_01259_)
);

NAND2_X1 _06268_ (
  .A1(_01258_),
  .A2(_01259_),
  .ZN(_00093_)
);

NAND2_X1 _06269_ (
  .A1(_01248_),
  .A2(\sresult[6][10] ),
  .ZN(_01260_)
);

NAND2_X1 _06270_ (
  .A1(_01237_),
  .A2(din_65[10]),
  .ZN(_01261_)
);

NAND2_X1 _06271_ (
  .A1(_01260_),
  .A2(_01261_),
  .ZN(_01262_)
);

NAND2_X1 _06272_ (
  .A1(_01262_),
  .A2(_01240_),
  .ZN(_01263_)
);

NAND2_X1 _06273_ (
  .A1(_01253_),
  .A2(\sresult[7][10] ),
  .ZN(_01264_)
);

NAND2_X1 _06274_ (
  .A1(_01263_),
  .A2(_01264_),
  .ZN(_00094_)
);

NAND2_X1 _06275_ (
  .A1(_01248_),
  .A2(\sresult[6][11] ),
  .ZN(_01265_)
);

NAND2_X1 _06276_ (
  .A1(_01237_),
  .A2(din_65[11]),
  .ZN(_01266_)
);

NAND2_X1 _06277_ (
  .A1(_01265_),
  .A2(_01266_),
  .ZN(_01267_)
);

NAND2_X1 _06278_ (
  .A1(_01267_),
  .A2(_01240_),
  .ZN(_01268_)
);

NAND2_X1 _06279_ (
  .A1(_01253_),
  .A2(\sresult[7][11] ),
  .ZN(_01269_)
);

NAND2_X1 _06280_ (
  .A1(_01268_),
  .A2(_01269_),
  .ZN(_00095_)
);

NAND2_X1 _06281_ (
  .A1(_01248_),
  .A2(\sresult[7][0] ),
  .ZN(_01270_)
);

NAND2_X1 _06282_ (
  .A1(_01237_),
  .A2(din_56[0]),
  .ZN(_01271_)
);

NAND2_X1 _06283_ (
  .A1(_01270_),
  .A2(_01271_),
  .ZN(_01272_)
);

NAND2_X1 _06284_ (
  .A1(_01272_),
  .A2(_01240_),
  .ZN(_01273_)
);

NAND2_X1 _06285_ (
  .A1(_01253_),
  .A2(\sresult[8][0] ),
  .ZN(_01274_)
);

NAND2_X1 _06286_ (
  .A1(_01273_),
  .A2(_01274_),
  .ZN(_00096_)
);

NAND2_X1 _06287_ (
  .A1(_01248_),
  .A2(\sresult[7][1] ),
  .ZN(_01275_)
);

NAND2_X1 _06288_ (
  .A1(_01237_),
  .A2(din_56[1]),
  .ZN(_01276_)
);

NAND2_X1 _06289_ (
  .A1(_01275_),
  .A2(_01276_),
  .ZN(_01277_)
);

NAND2_X1 _06290_ (
  .A1(_01277_),
  .A2(_01240_),
  .ZN(_01278_)
);

NAND2_X1 _06291_ (
  .A1(_01253_),
  .A2(\sresult[8][1] ),
  .ZN(_01279_)
);

NAND2_X1 _06292_ (
  .A1(_01278_),
  .A2(_01279_),
  .ZN(_00097_)
);

NAND2_X1 _06293_ (
  .A1(_01248_),
  .A2(\sresult[7][2] ),
  .ZN(_01280_)
);

NAND2_X1 _06294_ (
  .A1(_01237_),
  .A2(din_56[2]),
  .ZN(_01281_)
);

NAND2_X1 _06295_ (
  .A1(_01280_),
  .A2(_01281_),
  .ZN(_01282_)
);

NAND2_X1 _06296_ (
  .A1(_01282_),
  .A2(_01240_),
  .ZN(_01283_)
);

NAND2_X1 _06297_ (
  .A1(_01253_),
  .A2(\sresult[8][2] ),
  .ZN(_01284_)
);

NAND2_X1 _06298_ (
  .A1(_01283_),
  .A2(_01284_),
  .ZN(_00098_)
);

NAND2_X1 _06299_ (
  .A1(_01248_),
  .A2(\sresult[7][3] ),
  .ZN(_01285_)
);

NAND2_X1 _06300_ (
  .A1(_01237_),
  .A2(din_56[3]),
  .ZN(_01286_)
);

NAND2_X1 _06301_ (
  .A1(_01285_),
  .A2(_01286_),
  .ZN(_01287_)
);

NAND2_X1 _06302_ (
  .A1(_01287_),
  .A2(_01240_),
  .ZN(_01288_)
);

NAND2_X1 _06303_ (
  .A1(_01253_),
  .A2(\sresult[8][3] ),
  .ZN(_01289_)
);

NAND2_X1 _06304_ (
  .A1(_01288_),
  .A2(_01289_),
  .ZN(_00099_)
);

NAND2_X1 _06305_ (
  .A1(_01248_),
  .A2(\sresult[7][4] ),
  .ZN(_01290_)
);

BUF_X4 _06306_ (
  .A(_01019_),
  .Z(_01291_)
);

NAND2_X1 _06307_ (
  .A1(_01291_),
  .A2(din_56[4]),
  .ZN(_01292_)
);

NAND2_X1 _06308_ (
  .A1(_01290_),
  .A2(_01292_),
  .ZN(_01293_)
);

BUF_X2 _06309_ (
  .A(_00912_),
  .Z(_01294_)
);

NAND2_X1 _06310_ (
  .A1(_01293_),
  .A2(_01294_),
  .ZN(_01295_)
);

NAND2_X1 _06311_ (
  .A1(_01253_),
  .A2(\sresult[8][4] ),
  .ZN(_01296_)
);

NAND2_X1 _06312_ (
  .A1(_01295_),
  .A2(_01296_),
  .ZN(_00100_)
);

NAND2_X1 _06313_ (
  .A1(_01248_),
  .A2(\sresult[7][5] ),
  .ZN(_01297_)
);

NAND2_X1 _06314_ (
  .A1(_01291_),
  .A2(din_56[5]),
  .ZN(_01298_)
);

NAND2_X1 _06315_ (
  .A1(_01297_),
  .A2(_01298_),
  .ZN(_01299_)
);

NAND2_X1 _06316_ (
  .A1(_01299_),
  .A2(_01294_),
  .ZN(_01300_)
);

NAND2_X1 _06317_ (
  .A1(_01253_),
  .A2(\sresult[8][5] ),
  .ZN(_01301_)
);

NAND2_X1 _06318_ (
  .A1(_01300_),
  .A2(_01301_),
  .ZN(_00101_)
);

BUF_X4 _06319_ (
  .A(_00975_),
  .Z(_01302_)
);

NAND2_X1 _06320_ (
  .A1(_01302_),
  .A2(\sresult[7][6] ),
  .ZN(_01303_)
);

NAND2_X1 _06321_ (
  .A1(_01291_),
  .A2(din_56[6]),
  .ZN(_01304_)
);

NAND2_X1 _06322_ (
  .A1(_01303_),
  .A2(_01304_),
  .ZN(_01305_)
);

NAND2_X1 _06323_ (
  .A1(_01305_),
  .A2(_01294_),
  .ZN(_01306_)
);

CLKBUF_X2 _06324_ (
  .A(_01036_),
  .Z(_01307_)
);

NAND2_X1 _06325_ (
  .A1(_01307_),
  .A2(\sresult[8][6] ),
  .ZN(_01308_)
);

NAND2_X1 _06326_ (
  .A1(_01306_),
  .A2(_01308_),
  .ZN(_00102_)
);

NAND2_X1 _06327_ (
  .A1(_01302_),
  .A2(\sresult[7][7] ),
  .ZN(_01309_)
);

NAND2_X1 _06328_ (
  .A1(_01291_),
  .A2(din_56[7]),
  .ZN(_01310_)
);

NAND2_X1 _06329_ (
  .A1(_01309_),
  .A2(_01310_),
  .ZN(_01311_)
);

NAND2_X1 _06330_ (
  .A1(_01311_),
  .A2(_01294_),
  .ZN(_01312_)
);

NAND2_X1 _06331_ (
  .A1(_01307_),
  .A2(\sresult[8][7] ),
  .ZN(_01313_)
);

NAND2_X1 _06332_ (
  .A1(_01312_),
  .A2(_01313_),
  .ZN(_00103_)
);

NAND2_X1 _06333_ (
  .A1(_01302_),
  .A2(\sresult[7][8] ),
  .ZN(_01314_)
);

NAND2_X1 _06334_ (
  .A1(_01291_),
  .A2(din_56[8]),
  .ZN(_01315_)
);

NAND2_X1 _06335_ (
  .A1(_01314_),
  .A2(_01315_),
  .ZN(_01316_)
);

NAND2_X1 _06336_ (
  .A1(_01316_),
  .A2(_01294_),
  .ZN(_01317_)
);

NAND2_X1 _06337_ (
  .A1(_01307_),
  .A2(\sresult[8][8] ),
  .ZN(_01318_)
);

NAND2_X1 _06338_ (
  .A1(_01317_),
  .A2(_01318_),
  .ZN(_00104_)
);

NAND2_X1 _06339_ (
  .A1(_01302_),
  .A2(\sresult[7][9] ),
  .ZN(_01319_)
);

NAND2_X1 _06340_ (
  .A1(_01291_),
  .A2(din_56[9]),
  .ZN(_01320_)
);

NAND2_X1 _06341_ (
  .A1(_01319_),
  .A2(_01320_),
  .ZN(_01321_)
);

NAND2_X1 _06342_ (
  .A1(_01321_),
  .A2(_01294_),
  .ZN(_01322_)
);

NAND2_X1 _06343_ (
  .A1(_01307_),
  .A2(\sresult[8][9] ),
  .ZN(_01323_)
);

NAND2_X1 _06344_ (
  .A1(_01322_),
  .A2(_01323_),
  .ZN(_00105_)
);

NAND2_X1 _06345_ (
  .A1(_01302_),
  .A2(\sresult[7][10] ),
  .ZN(_01324_)
);

NAND2_X1 _06346_ (
  .A1(_01291_),
  .A2(din_56[10]),
  .ZN(_01325_)
);

NAND2_X1 _06347_ (
  .A1(_01324_),
  .A2(_01325_),
  .ZN(_01326_)
);

NAND2_X1 _06348_ (
  .A1(_01326_),
  .A2(_01294_),
  .ZN(_01327_)
);

NAND2_X1 _06349_ (
  .A1(_01307_),
  .A2(\sresult[8][10] ),
  .ZN(_01328_)
);

NAND2_X1 _06350_ (
  .A1(_01327_),
  .A2(_01328_),
  .ZN(_00106_)
);

NAND2_X1 _06351_ (
  .A1(_01302_),
  .A2(\sresult[7][11] ),
  .ZN(_01329_)
);

NAND2_X1 _06352_ (
  .A1(_01291_),
  .A2(din_56[11]),
  .ZN(_01330_)
);

NAND2_X1 _06353_ (
  .A1(_01329_),
  .A2(_01330_),
  .ZN(_01331_)
);

NAND2_X1 _06354_ (
  .A1(_01331_),
  .A2(_01294_),
  .ZN(_01332_)
);

NAND2_X1 _06355_ (
  .A1(_01307_),
  .A2(\sresult[8][11] ),
  .ZN(_01333_)
);

NAND2_X1 _06356_ (
  .A1(_01332_),
  .A2(_01333_),
  .ZN(_00107_)
);

NAND2_X1 _06357_ (
  .A1(_01302_),
  .A2(\sresult[8][0] ),
  .ZN(_01334_)
);

NAND2_X1 _06358_ (
  .A1(_01291_),
  .A2(din_47[0]),
  .ZN(_01335_)
);

NAND2_X1 _06359_ (
  .A1(_01334_),
  .A2(_01335_),
  .ZN(_01336_)
);

NAND2_X1 _06360_ (
  .A1(_01336_),
  .A2(_01294_),
  .ZN(_01337_)
);

NAND2_X1 _06361_ (
  .A1(_01307_),
  .A2(\sresult[9][0] ),
  .ZN(_01338_)
);

NAND2_X1 _06362_ (
  .A1(_01337_),
  .A2(_01338_),
  .ZN(_00108_)
);

NAND2_X1 _06363_ (
  .A1(_01302_),
  .A2(\sresult[8][1] ),
  .ZN(_01339_)
);

NAND2_X1 _06364_ (
  .A1(_01291_),
  .A2(din_47[1]),
  .ZN(_01340_)
);

NAND2_X1 _06365_ (
  .A1(_01339_),
  .A2(_01340_),
  .ZN(_01341_)
);

NAND2_X1 _06366_ (
  .A1(_01341_),
  .A2(_01294_),
  .ZN(_01342_)
);

NAND2_X1 _06367_ (
  .A1(_01307_),
  .A2(\sresult[9][1] ),
  .ZN(_01343_)
);

NAND2_X1 _06368_ (
  .A1(_01342_),
  .A2(_01343_),
  .ZN(_00109_)
);

NAND2_X1 _06369_ (
  .A1(_01302_),
  .A2(\sresult[8][2] ),
  .ZN(_01344_)
);

BUF_X4 _06370_ (
  .A(_01019_),
  .Z(_01345_)
);

NAND2_X1 _06371_ (
  .A1(_01345_),
  .A2(din_47[2]),
  .ZN(_01346_)
);

NAND2_X1 _06372_ (
  .A1(_01344_),
  .A2(_01346_),
  .ZN(_01347_)
);

BUF_X2 _06373_ (
  .A(_00912_),
  .Z(_01348_)
);

NAND2_X1 _06374_ (
  .A1(_01347_),
  .A2(_01348_),
  .ZN(_01349_)
);

NAND2_X1 _06375_ (
  .A1(_01307_),
  .A2(\sresult[9][2] ),
  .ZN(_01350_)
);

NAND2_X1 _06376_ (
  .A1(_01349_),
  .A2(_01350_),
  .ZN(_00110_)
);

NAND2_X1 _06377_ (
  .A1(_01302_),
  .A2(\sresult[8][3] ),
  .ZN(_01351_)
);

NAND2_X1 _06378_ (
  .A1(_01345_),
  .A2(din_47[3]),
  .ZN(_01352_)
);

NAND2_X1 _06379_ (
  .A1(_01351_),
  .A2(_01352_),
  .ZN(_01353_)
);

NAND2_X1 _06380_ (
  .A1(_01353_),
  .A2(_01348_),
  .ZN(_01354_)
);

NAND2_X1 _06381_ (
  .A1(_01307_),
  .A2(\sresult[9][3] ),
  .ZN(_01355_)
);

NAND2_X1 _06382_ (
  .A1(_01354_),
  .A2(_01355_),
  .ZN(_00111_)
);

BUF_X4 _06383_ (
  .A(_00975_),
  .Z(_01356_)
);

NAND2_X1 _06384_ (
  .A1(_01356_),
  .A2(\sresult[8][4] ),
  .ZN(_01357_)
);

NAND2_X1 _06385_ (
  .A1(_01345_),
  .A2(din_47[4]),
  .ZN(_01358_)
);

NAND2_X1 _06386_ (
  .A1(_01357_),
  .A2(_01358_),
  .ZN(_01359_)
);

NAND2_X1 _06387_ (
  .A1(_01359_),
  .A2(_01348_),
  .ZN(_01360_)
);

CLKBUF_X2 _06388_ (
  .A(_01036_),
  .Z(_01361_)
);

NAND2_X1 _06389_ (
  .A1(_01361_),
  .A2(\sresult[9][4] ),
  .ZN(_01362_)
);

NAND2_X1 _06390_ (
  .A1(_01360_),
  .A2(_01362_),
  .ZN(_00112_)
);

NAND2_X1 _06391_ (
  .A1(_01356_),
  .A2(\sresult[8][5] ),
  .ZN(_01363_)
);

NAND2_X1 _06392_ (
  .A1(_01345_),
  .A2(din_47[5]),
  .ZN(_01364_)
);

NAND2_X1 _06393_ (
  .A1(_01363_),
  .A2(_01364_),
  .ZN(_01365_)
);

NAND2_X1 _06394_ (
  .A1(_01365_),
  .A2(_01348_),
  .ZN(_01366_)
);

NAND2_X1 _06395_ (
  .A1(_01361_),
  .A2(\sresult[9][5] ),
  .ZN(_01367_)
);

NAND2_X1 _06396_ (
  .A1(_01366_),
  .A2(_01367_),
  .ZN(_00113_)
);

NAND2_X1 _06397_ (
  .A1(_01356_),
  .A2(\sresult[8][6] ),
  .ZN(_01368_)
);

NAND2_X1 _06398_ (
  .A1(_01345_),
  .A2(din_47[6]),
  .ZN(_01369_)
);

NAND2_X1 _06399_ (
  .A1(_01368_),
  .A2(_01369_),
  .ZN(_01370_)
);

NAND2_X1 _06400_ (
  .A1(_01370_),
  .A2(_01348_),
  .ZN(_01371_)
);

NAND2_X1 _06401_ (
  .A1(_01361_),
  .A2(\sresult[9][6] ),
  .ZN(_01372_)
);

NAND2_X1 _06402_ (
  .A1(_01371_),
  .A2(_01372_),
  .ZN(_00114_)
);

NAND2_X1 _06403_ (
  .A1(_01356_),
  .A2(\sresult[8][7] ),
  .ZN(_01373_)
);

NAND2_X1 _06404_ (
  .A1(_01345_),
  .A2(din_47[7]),
  .ZN(_01374_)
);

NAND2_X1 _06405_ (
  .A1(_01373_),
  .A2(_01374_),
  .ZN(_01375_)
);

NAND2_X1 _06406_ (
  .A1(_01375_),
  .A2(_01348_),
  .ZN(_01376_)
);

NAND2_X1 _06407_ (
  .A1(_01361_),
  .A2(\sresult[9][7] ),
  .ZN(_01377_)
);

NAND2_X1 _06408_ (
  .A1(_01376_),
  .A2(_01377_),
  .ZN(_00115_)
);

NAND2_X1 _06409_ (
  .A1(_01356_),
  .A2(\sresult[8][8] ),
  .ZN(_01378_)
);

NAND2_X1 _06410_ (
  .A1(_01345_),
  .A2(din_47[8]),
  .ZN(_01379_)
);

NAND2_X1 _06411_ (
  .A1(_01378_),
  .A2(_01379_),
  .ZN(_01380_)
);

NAND2_X1 _06412_ (
  .A1(_01380_),
  .A2(_01348_),
  .ZN(_01381_)
);

NAND2_X1 _06413_ (
  .A1(_01361_),
  .A2(\sresult[9][8] ),
  .ZN(_01382_)
);

NAND2_X1 _06414_ (
  .A1(_01381_),
  .A2(_01382_),
  .ZN(_00116_)
);

NAND2_X1 _06415_ (
  .A1(_01356_),
  .A2(\sresult[8][9] ),
  .ZN(_01383_)
);

NAND2_X1 _06416_ (
  .A1(_01345_),
  .A2(din_47[9]),
  .ZN(_01384_)
);

NAND2_X1 _06417_ (
  .A1(_01383_),
  .A2(_01384_),
  .ZN(_01385_)
);

NAND2_X1 _06418_ (
  .A1(_01385_),
  .A2(_01348_),
  .ZN(_01386_)
);

NAND2_X1 _06419_ (
  .A1(_01361_),
  .A2(\sresult[9][9] ),
  .ZN(_01387_)
);

NAND2_X1 _06420_ (
  .A1(_01386_),
  .A2(_01387_),
  .ZN(_00117_)
);

NAND2_X1 _06421_ (
  .A1(_01356_),
  .A2(\sresult[8][10] ),
  .ZN(_01388_)
);

NAND2_X1 _06422_ (
  .A1(_01345_),
  .A2(din_47[10]),
  .ZN(_01389_)
);

NAND2_X1 _06423_ (
  .A1(_01388_),
  .A2(_01389_),
  .ZN(_01390_)
);

NAND2_X1 _06424_ (
  .A1(_01390_),
  .A2(_01348_),
  .ZN(_01391_)
);

NAND2_X1 _06425_ (
  .A1(_01361_),
  .A2(\sresult[9][10] ),
  .ZN(_01392_)
);

NAND2_X1 _06426_ (
  .A1(_01391_),
  .A2(_01392_),
  .ZN(_00118_)
);

NAND2_X1 _06427_ (
  .A1(_01356_),
  .A2(\sresult[8][11] ),
  .ZN(_01393_)
);

NAND2_X1 _06428_ (
  .A1(_01345_),
  .A2(din_47[11]),
  .ZN(_01394_)
);

NAND2_X1 _06429_ (
  .A1(_01393_),
  .A2(_01394_),
  .ZN(_01395_)
);

NAND2_X1 _06430_ (
  .A1(_01395_),
  .A2(_01348_),
  .ZN(_01396_)
);

NAND2_X1 _06431_ (
  .A1(_01361_),
  .A2(\sresult[9][11] ),
  .ZN(_01397_)
);

NAND2_X1 _06432_ (
  .A1(_01396_),
  .A2(_01397_),
  .ZN(_00119_)
);

NAND2_X1 _06433_ (
  .A1(_01356_),
  .A2(\sresult[9][0] ),
  .ZN(_01398_)
);

BUF_X4 _06434_ (
  .A(_01019_),
  .Z(_01399_)
);

NAND2_X1 _06435_ (
  .A1(_01399_),
  .A2(din_37[0]),
  .ZN(_01400_)
);

NAND2_X1 _06436_ (
  .A1(_01398_),
  .A2(_01400_),
  .ZN(_01401_)
);

BUF_X2 _06437_ (
  .A(_00912_),
  .Z(_01402_)
);

NAND2_X1 _06438_ (
  .A1(_01401_),
  .A2(_01402_),
  .ZN(_01403_)
);

NAND2_X1 _06439_ (
  .A1(_01361_),
  .A2(\sresult[10][0] ),
  .ZN(_01404_)
);

NAND2_X1 _06440_ (
  .A1(_01403_),
  .A2(_01404_),
  .ZN(_00120_)
);

NAND2_X1 _06441_ (
  .A1(_01356_),
  .A2(\sresult[9][1] ),
  .ZN(_01405_)
);

NAND2_X1 _06442_ (
  .A1(_01399_),
  .A2(din_37[1]),
  .ZN(_01406_)
);

NAND2_X1 _06443_ (
  .A1(_01405_),
  .A2(_01406_),
  .ZN(_01407_)
);

NAND2_X1 _06444_ (
  .A1(_01407_),
  .A2(_01402_),
  .ZN(_01408_)
);

NAND2_X1 _06445_ (
  .A1(_01361_),
  .A2(\sresult[10][1] ),
  .ZN(_01409_)
);

NAND2_X1 _06446_ (
  .A1(_01408_),
  .A2(_01409_),
  .ZN(_00121_)
);

BUF_X4 _06447_ (
  .A(_00975_),
  .Z(_01410_)
);

NAND2_X1 _06448_ (
  .A1(_01410_),
  .A2(\sresult[9][2] ),
  .ZN(_01411_)
);

NAND2_X1 _06449_ (
  .A1(_01399_),
  .A2(din_37[2]),
  .ZN(_01412_)
);

NAND2_X1 _06450_ (
  .A1(_01411_),
  .A2(_01412_),
  .ZN(_01413_)
);

NAND2_X1 _06451_ (
  .A1(_01413_),
  .A2(_01402_),
  .ZN(_01414_)
);

CLKBUF_X2 _06452_ (
  .A(_01036_),
  .Z(_01415_)
);

NAND2_X1 _06453_ (
  .A1(_01415_),
  .A2(\sresult[10][2] ),
  .ZN(_01416_)
);

NAND2_X1 _06454_ (
  .A1(_01414_),
  .A2(_01416_),
  .ZN(_00122_)
);

NAND2_X1 _06455_ (
  .A1(_01410_),
  .A2(\sresult[9][3] ),
  .ZN(_01417_)
);

NAND2_X1 _06456_ (
  .A1(_01399_),
  .A2(din_37[3]),
  .ZN(_01418_)
);

NAND2_X1 _06457_ (
  .A1(_01417_),
  .A2(_01418_),
  .ZN(_01419_)
);

NAND2_X1 _06458_ (
  .A1(_01419_),
  .A2(_01402_),
  .ZN(_01420_)
);

NAND2_X1 _06459_ (
  .A1(_01415_),
  .A2(\sresult[10][3] ),
  .ZN(_01421_)
);

NAND2_X1 _06460_ (
  .A1(_01420_),
  .A2(_01421_),
  .ZN(_00123_)
);

NAND2_X1 _06461_ (
  .A1(_01410_),
  .A2(\sresult[9][4] ),
  .ZN(_01422_)
);

NAND2_X1 _06462_ (
  .A1(_01399_),
  .A2(din_37[4]),
  .ZN(_01423_)
);

NAND2_X1 _06463_ (
  .A1(_01422_),
  .A2(_01423_),
  .ZN(_01424_)
);

NAND2_X1 _06464_ (
  .A1(_01424_),
  .A2(_01402_),
  .ZN(_01425_)
);

NAND2_X1 _06465_ (
  .A1(_01415_),
  .A2(\sresult[10][4] ),
  .ZN(_01426_)
);

NAND2_X1 _06466_ (
  .A1(_01425_),
  .A2(_01426_),
  .ZN(_00124_)
);

NAND2_X1 _06467_ (
  .A1(_01410_),
  .A2(\sresult[9][5] ),
  .ZN(_01427_)
);

NAND2_X1 _06468_ (
  .A1(_01399_),
  .A2(din_37[5]),
  .ZN(_01428_)
);

NAND2_X1 _06469_ (
  .A1(_01427_),
  .A2(_01428_),
  .ZN(_01429_)
);

NAND2_X1 _06470_ (
  .A1(_01429_),
  .A2(_01402_),
  .ZN(_01430_)
);

NAND2_X1 _06471_ (
  .A1(_01415_),
  .A2(\sresult[10][5] ),
  .ZN(_01431_)
);

NAND2_X1 _06472_ (
  .A1(_01430_),
  .A2(_01431_),
  .ZN(_00125_)
);

NAND2_X1 _06473_ (
  .A1(_01410_),
  .A2(\sresult[9][6] ),
  .ZN(_01432_)
);

NAND2_X1 _06474_ (
  .A1(_01399_),
  .A2(din_37[6]),
  .ZN(_01433_)
);

NAND2_X1 _06475_ (
  .A1(_01432_),
  .A2(_01433_),
  .ZN(_01434_)
);

NAND2_X1 _06476_ (
  .A1(_01434_),
  .A2(_01402_),
  .ZN(_01435_)
);

NAND2_X1 _06477_ (
  .A1(_01415_),
  .A2(\sresult[10][6] ),
  .ZN(_01436_)
);

NAND2_X1 _06478_ (
  .A1(_01435_),
  .A2(_01436_),
  .ZN(_00126_)
);

NAND2_X1 _06479_ (
  .A1(_01410_),
  .A2(\sresult[9][7] ),
  .ZN(_01437_)
);

NAND2_X1 _06480_ (
  .A1(_01399_),
  .A2(din_37[7]),
  .ZN(_01438_)
);

NAND2_X1 _06481_ (
  .A1(_01437_),
  .A2(_01438_),
  .ZN(_01439_)
);

NAND2_X1 _06482_ (
  .A1(_01439_),
  .A2(_01402_),
  .ZN(_01440_)
);

NAND2_X1 _06483_ (
  .A1(_01415_),
  .A2(\sresult[10][7] ),
  .ZN(_01441_)
);

NAND2_X1 _06484_ (
  .A1(_01440_),
  .A2(_01441_),
  .ZN(_00127_)
);

NAND2_X1 _06485_ (
  .A1(_01410_),
  .A2(\sresult[9][8] ),
  .ZN(_01442_)
);

NAND2_X1 _06486_ (
  .A1(_01399_),
  .A2(din_37[8]),
  .ZN(_01443_)
);

NAND2_X1 _06487_ (
  .A1(_01442_),
  .A2(_01443_),
  .ZN(_01444_)
);

NAND2_X1 _06488_ (
  .A1(_01444_),
  .A2(_01402_),
  .ZN(_01445_)
);

NAND2_X1 _06489_ (
  .A1(_01415_),
  .A2(\sresult[10][8] ),
  .ZN(_01446_)
);

NAND2_X1 _06490_ (
  .A1(_01445_),
  .A2(_01446_),
  .ZN(_00128_)
);

NAND2_X1 _06491_ (
  .A1(_01410_),
  .A2(\sresult[9][9] ),
  .ZN(_01447_)
);

NAND2_X1 _06492_ (
  .A1(_01399_),
  .A2(din_37[9]),
  .ZN(_01448_)
);

NAND2_X1 _06493_ (
  .A1(_01447_),
  .A2(_01448_),
  .ZN(_01449_)
);

NAND2_X1 _06494_ (
  .A1(_01449_),
  .A2(_01402_),
  .ZN(_01450_)
);

NAND2_X1 _06495_ (
  .A1(_01415_),
  .A2(\sresult[10][9] ),
  .ZN(_01451_)
);

NAND2_X1 _06496_ (
  .A1(_01450_),
  .A2(_01451_),
  .ZN(_00129_)
);

NAND2_X1 _06497_ (
  .A1(_01410_),
  .A2(\sresult[9][10] ),
  .ZN(_01452_)
);

BUF_X4 _06498_ (
  .A(_01019_),
  .Z(_01453_)
);

NAND2_X1 _06499_ (
  .A1(_01453_),
  .A2(din_37[10]),
  .ZN(_01454_)
);

NAND2_X1 _06500_ (
  .A1(_01452_),
  .A2(_01454_),
  .ZN(_01455_)
);

BUF_X4 _06501_ (
  .A(_00911_),
  .Z(_01456_)
);

BUF_X2 _06502_ (
  .A(_01456_),
  .Z(_01457_)
);

NAND2_X1 _06503_ (
  .A1(_01455_),
  .A2(_01457_),
  .ZN(_01458_)
);

NAND2_X1 _06504_ (
  .A1(_01415_),
  .A2(\sresult[10][10] ),
  .ZN(_01459_)
);

NAND2_X1 _06505_ (
  .A1(_01458_),
  .A2(_01459_),
  .ZN(_00130_)
);

NAND2_X1 _06506_ (
  .A1(_01410_),
  .A2(\sresult[9][11] ),
  .ZN(_01460_)
);

NAND2_X1 _06507_ (
  .A1(_01453_),
  .A2(din_37[11]),
  .ZN(_01461_)
);

NAND2_X1 _06508_ (
  .A1(_01460_),
  .A2(_01461_),
  .ZN(_01462_)
);

NAND2_X1 _06509_ (
  .A1(_01462_),
  .A2(_01457_),
  .ZN(_01463_)
);

NAND2_X1 _06510_ (
  .A1(_01415_),
  .A2(\sresult[10][11] ),
  .ZN(_01464_)
);

NAND2_X1 _06511_ (
  .A1(_01463_),
  .A2(_01464_),
  .ZN(_00131_)
);

BUF_X4 _06512_ (
  .A(_00975_),
  .Z(_01465_)
);

NAND2_X1 _06513_ (
  .A1(_01465_),
  .A2(\sresult[10][0] ),
  .ZN(_01466_)
);

NAND2_X1 _06514_ (
  .A1(_01453_),
  .A2(din_46[0]),
  .ZN(_01467_)
);

NAND2_X1 _06515_ (
  .A1(_01466_),
  .A2(_01467_),
  .ZN(_01468_)
);

NAND2_X1 _06516_ (
  .A1(_01468_),
  .A2(_01457_),
  .ZN(_01469_)
);

CLKBUF_X2 _06517_ (
  .A(_01036_),
  .Z(_01470_)
);

NAND2_X1 _06518_ (
  .A1(_01470_),
  .A2(\sresult[11][0] ),
  .ZN(_01471_)
);

NAND2_X1 _06519_ (
  .A1(_01469_),
  .A2(_01471_),
  .ZN(_00132_)
);

NAND2_X1 _06520_ (
  .A1(_01465_),
  .A2(\sresult[10][1] ),
  .ZN(_01472_)
);

NAND2_X1 _06521_ (
  .A1(_01453_),
  .A2(din_46[1]),
  .ZN(_01473_)
);

NAND2_X1 _06522_ (
  .A1(_01472_),
  .A2(_01473_),
  .ZN(_01474_)
);

NAND2_X1 _06523_ (
  .A1(_01474_),
  .A2(_01457_),
  .ZN(_01475_)
);

NAND2_X1 _06524_ (
  .A1(_01470_),
  .A2(\sresult[11][1] ),
  .ZN(_01476_)
);

NAND2_X1 _06525_ (
  .A1(_01475_),
  .A2(_01476_),
  .ZN(_00133_)
);

NAND2_X1 _06526_ (
  .A1(_01465_),
  .A2(\sresult[10][2] ),
  .ZN(_01477_)
);

NAND2_X1 _06527_ (
  .A1(_01453_),
  .A2(din_46[2]),
  .ZN(_01478_)
);

NAND2_X1 _06528_ (
  .A1(_01477_),
  .A2(_01478_),
  .ZN(_01479_)
);

NAND2_X1 _06529_ (
  .A1(_01479_),
  .A2(_01457_),
  .ZN(_01480_)
);

NAND2_X1 _06530_ (
  .A1(_01470_),
  .A2(\sresult[11][2] ),
  .ZN(_01481_)
);

NAND2_X1 _06531_ (
  .A1(_01480_),
  .A2(_01481_),
  .ZN(_00134_)
);

NAND2_X1 _06532_ (
  .A1(_01465_),
  .A2(\sresult[10][3] ),
  .ZN(_01482_)
);

NAND2_X1 _06533_ (
  .A1(_01453_),
  .A2(din_46[3]),
  .ZN(_01483_)
);

NAND2_X1 _06534_ (
  .A1(_01482_),
  .A2(_01483_),
  .ZN(_01484_)
);

NAND2_X1 _06535_ (
  .A1(_01484_),
  .A2(_01457_),
  .ZN(_01485_)
);

NAND2_X1 _06536_ (
  .A1(_01470_),
  .A2(\sresult[11][3] ),
  .ZN(_01486_)
);

NAND2_X1 _06537_ (
  .A1(_01485_),
  .A2(_01486_),
  .ZN(_00135_)
);

NAND2_X1 _06538_ (
  .A1(_01465_),
  .A2(\sresult[10][4] ),
  .ZN(_01487_)
);

NAND2_X1 _06539_ (
  .A1(_01453_),
  .A2(din_46[4]),
  .ZN(_01488_)
);

NAND2_X1 _06540_ (
  .A1(_01487_),
  .A2(_01488_),
  .ZN(_01489_)
);

NAND2_X1 _06541_ (
  .A1(_01489_),
  .A2(_01457_),
  .ZN(_01490_)
);

NAND2_X1 _06542_ (
  .A1(_01470_),
  .A2(\sresult[11][4] ),
  .ZN(_01491_)
);

NAND2_X1 _06543_ (
  .A1(_01490_),
  .A2(_01491_),
  .ZN(_00136_)
);

NAND2_X1 _06544_ (
  .A1(_01465_),
  .A2(\sresult[10][5] ),
  .ZN(_01492_)
);

NAND2_X1 _06545_ (
  .A1(_01453_),
  .A2(din_46[5]),
  .ZN(_01493_)
);

NAND2_X1 _06546_ (
  .A1(_01492_),
  .A2(_01493_),
  .ZN(_01494_)
);

NAND2_X1 _06547_ (
  .A1(_01494_),
  .A2(_01457_),
  .ZN(_01495_)
);

NAND2_X1 _06548_ (
  .A1(_01470_),
  .A2(\sresult[11][5] ),
  .ZN(_01496_)
);

NAND2_X1 _06549_ (
  .A1(_01495_),
  .A2(_01496_),
  .ZN(_00137_)
);

NAND2_X1 _06550_ (
  .A1(_01465_),
  .A2(\sresult[10][6] ),
  .ZN(_01497_)
);

NAND2_X1 _06551_ (
  .A1(_01453_),
  .A2(din_46[6]),
  .ZN(_01498_)
);

NAND2_X1 _06552_ (
  .A1(_01497_),
  .A2(_01498_),
  .ZN(_01499_)
);

NAND2_X1 _06553_ (
  .A1(_01499_),
  .A2(_01457_),
  .ZN(_01500_)
);

NAND2_X1 _06554_ (
  .A1(_01470_),
  .A2(\sresult[11][6] ),
  .ZN(_01501_)
);

NAND2_X1 _06555_ (
  .A1(_01500_),
  .A2(_01501_),
  .ZN(_00138_)
);

NAND2_X1 _06556_ (
  .A1(_01465_),
  .A2(\sresult[10][7] ),
  .ZN(_01502_)
);

NAND2_X1 _06557_ (
  .A1(_01453_),
  .A2(din_46[7]),
  .ZN(_01503_)
);

NAND2_X1 _06558_ (
  .A1(_01502_),
  .A2(_01503_),
  .ZN(_01504_)
);

NAND2_X1 _06559_ (
  .A1(_01504_),
  .A2(_01457_),
  .ZN(_01505_)
);

NAND2_X1 _06560_ (
  .A1(_01470_),
  .A2(\sresult[11][7] ),
  .ZN(_01506_)
);

NAND2_X1 _06561_ (
  .A1(_01505_),
  .A2(_01506_),
  .ZN(_00139_)
);

NAND2_X1 _06562_ (
  .A1(_01465_),
  .A2(\sresult[10][8] ),
  .ZN(_01507_)
);

BUF_X4 _06563_ (
  .A(_01019_),
  .Z(_01508_)
);

NAND2_X1 _06564_ (
  .A1(_01508_),
  .A2(din_46[8]),
  .ZN(_01509_)
);

NAND2_X1 _06565_ (
  .A1(_01507_),
  .A2(_01509_),
  .ZN(_01510_)
);

BUF_X2 _06566_ (
  .A(_01456_),
  .Z(_01511_)
);

NAND2_X1 _06567_ (
  .A1(_01510_),
  .A2(_01511_),
  .ZN(_01512_)
);

NAND2_X1 _06568_ (
  .A1(_01470_),
  .A2(\sresult[11][8] ),
  .ZN(_01513_)
);

NAND2_X1 _06569_ (
  .A1(_01512_),
  .A2(_01513_),
  .ZN(_00140_)
);

NAND2_X1 _06570_ (
  .A1(_01465_),
  .A2(\sresult[10][9] ),
  .ZN(_01514_)
);

NAND2_X1 _06571_ (
  .A1(_01508_),
  .A2(din_46[9]),
  .ZN(_01515_)
);

NAND2_X1 _06572_ (
  .A1(_01514_),
  .A2(_01515_),
  .ZN(_01516_)
);

NAND2_X1 _06573_ (
  .A1(_01516_),
  .A2(_01511_),
  .ZN(_01517_)
);

NAND2_X1 _06574_ (
  .A1(_01470_),
  .A2(\sresult[11][9] ),
  .ZN(_01518_)
);

NAND2_X1 _06575_ (
  .A1(_01517_),
  .A2(_01518_),
  .ZN(_00141_)
);

BUF_X8 _06576_ (
  .A(_00799_),
  .Z(_01519_)
);

BUF_X4 _06577_ (
  .A(_01519_),
  .Z(_01520_)
);

NAND2_X1 _06578_ (
  .A1(_01520_),
  .A2(\sresult[10][10] ),
  .ZN(_01521_)
);

NAND2_X1 _06579_ (
  .A1(_01508_),
  .A2(din_46[10]),
  .ZN(_01522_)
);

NAND2_X1 _06580_ (
  .A1(_01521_),
  .A2(_01522_),
  .ZN(_01523_)
);

NAND2_X1 _06581_ (
  .A1(_01523_),
  .A2(_01511_),
  .ZN(_01524_)
);

CLKBUF_X2 _06582_ (
  .A(_01036_),
  .Z(_01525_)
);

NAND2_X1 _06583_ (
  .A1(_01525_),
  .A2(\sresult[11][10] ),
  .ZN(_01526_)
);

NAND2_X1 _06584_ (
  .A1(_01524_),
  .A2(_01526_),
  .ZN(_00142_)
);

NAND2_X1 _06585_ (
  .A1(_01520_),
  .A2(\sresult[10][11] ),
  .ZN(_01527_)
);

NAND2_X1 _06586_ (
  .A1(_01508_),
  .A2(din_46[11]),
  .ZN(_01528_)
);

NAND2_X1 _06587_ (
  .A1(_01527_),
  .A2(_01528_),
  .ZN(_01529_)
);

NAND2_X1 _06588_ (
  .A1(_01529_),
  .A2(_01511_),
  .ZN(_01530_)
);

NAND2_X1 _06589_ (
  .A1(_01525_),
  .A2(\sresult[11][11] ),
  .ZN(_01531_)
);

NAND2_X1 _06590_ (
  .A1(_01530_),
  .A2(_01531_),
  .ZN(_00143_)
);

NAND2_X1 _06591_ (
  .A1(_01520_),
  .A2(\sresult[11][0] ),
  .ZN(_01532_)
);

NAND2_X1 _06592_ (
  .A1(_01508_),
  .A2(din_55[0]),
  .ZN(_01533_)
);

NAND2_X1 _06593_ (
  .A1(_01532_),
  .A2(_01533_),
  .ZN(_01534_)
);

NAND2_X1 _06594_ (
  .A1(_01534_),
  .A2(_01511_),
  .ZN(_01535_)
);

NAND2_X1 _06595_ (
  .A1(_01525_),
  .A2(\sresult[12][0] ),
  .ZN(_01536_)
);

NAND2_X1 _06596_ (
  .A1(_01535_),
  .A2(_01536_),
  .ZN(_00144_)
);

NAND2_X1 _06597_ (
  .A1(_01520_),
  .A2(\sresult[11][1] ),
  .ZN(_01537_)
);

NAND2_X1 _06598_ (
  .A1(_01508_),
  .A2(din_55[1]),
  .ZN(_01538_)
);

NAND2_X1 _06599_ (
  .A1(_01537_),
  .A2(_01538_),
  .ZN(_01539_)
);

NAND2_X1 _06600_ (
  .A1(_01539_),
  .A2(_01511_),
  .ZN(_01540_)
);

NAND2_X1 _06601_ (
  .A1(_01525_),
  .A2(\sresult[12][1] ),
  .ZN(_01541_)
);

NAND2_X1 _06602_ (
  .A1(_01540_),
  .A2(_01541_),
  .ZN(_00145_)
);

NAND2_X1 _06603_ (
  .A1(_01520_),
  .A2(\sresult[11][2] ),
  .ZN(_01542_)
);

NAND2_X1 _06604_ (
  .A1(_01508_),
  .A2(din_55[2]),
  .ZN(_01543_)
);

NAND2_X1 _06605_ (
  .A1(_01542_),
  .A2(_01543_),
  .ZN(_01544_)
);

NAND2_X1 _06606_ (
  .A1(_01544_),
  .A2(_01511_),
  .ZN(_01545_)
);

NAND2_X1 _06607_ (
  .A1(_01525_),
  .A2(\sresult[12][2] ),
  .ZN(_01546_)
);

NAND2_X1 _06608_ (
  .A1(_01545_),
  .A2(_01546_),
  .ZN(_00146_)
);

NAND2_X1 _06609_ (
  .A1(_01520_),
  .A2(\sresult[11][3] ),
  .ZN(_01547_)
);

NAND2_X1 _06610_ (
  .A1(_01508_),
  .A2(din_55[3]),
  .ZN(_01548_)
);

NAND2_X1 _06611_ (
  .A1(_01547_),
  .A2(_01548_),
  .ZN(_01549_)
);

NAND2_X1 _06612_ (
  .A1(_01549_),
  .A2(_01511_),
  .ZN(_01550_)
);

NAND2_X1 _06613_ (
  .A1(_01525_),
  .A2(\sresult[12][3] ),
  .ZN(_01551_)
);

NAND2_X1 _06614_ (
  .A1(_01550_),
  .A2(_01551_),
  .ZN(_00147_)
);

NAND2_X1 _06615_ (
  .A1(_01520_),
  .A2(\sresult[11][4] ),
  .ZN(_01552_)
);

NAND2_X1 _06616_ (
  .A1(_01508_),
  .A2(din_55[4]),
  .ZN(_01553_)
);

NAND2_X1 _06617_ (
  .A1(_01552_),
  .A2(_01553_),
  .ZN(_01554_)
);

NAND2_X1 _06618_ (
  .A1(_01554_),
  .A2(_01511_),
  .ZN(_01555_)
);

NAND2_X1 _06619_ (
  .A1(_01525_),
  .A2(\sresult[12][4] ),
  .ZN(_01556_)
);

NAND2_X1 _06620_ (
  .A1(_01555_),
  .A2(_01556_),
  .ZN(_00148_)
);

NAND2_X1 _06621_ (
  .A1(_01520_),
  .A2(\sresult[11][5] ),
  .ZN(_01557_)
);

NAND2_X1 _06622_ (
  .A1(_01508_),
  .A2(din_55[5]),
  .ZN(_01558_)
);

NAND2_X1 _06623_ (
  .A1(_01557_),
  .A2(_01558_),
  .ZN(_01559_)
);

NAND2_X1 _06624_ (
  .A1(_01559_),
  .A2(_01511_),
  .ZN(_01560_)
);

NAND2_X1 _06625_ (
  .A1(_01525_),
  .A2(\sresult[12][5] ),
  .ZN(_01561_)
);

NAND2_X1 _06626_ (
  .A1(_01560_),
  .A2(_01561_),
  .ZN(_00149_)
);

NAND2_X1 _06627_ (
  .A1(_01520_),
  .A2(\sresult[11][6] ),
  .ZN(_01562_)
);

BUF_X8 _06628_ (
  .A(_00770_),
  .Z(_01563_)
);

BUF_X4 _06629_ (
  .A(_01563_),
  .Z(_01564_)
);

NAND2_X1 _06630_ (
  .A1(_01564_),
  .A2(din_55[6]),
  .ZN(_01565_)
);

NAND2_X1 _06631_ (
  .A1(_01562_),
  .A2(_01565_),
  .ZN(_01566_)
);

BUF_X2 _06632_ (
  .A(_01456_),
  .Z(_01567_)
);

NAND2_X1 _06633_ (
  .A1(_01566_),
  .A2(_01567_),
  .ZN(_01568_)
);

NAND2_X1 _06634_ (
  .A1(_01525_),
  .A2(\sresult[12][6] ),
  .ZN(_01569_)
);

NAND2_X1 _06635_ (
  .A1(_01568_),
  .A2(_01569_),
  .ZN(_00150_)
);

NAND2_X1 _06636_ (
  .A1(_01520_),
  .A2(\sresult[11][7] ),
  .ZN(_01570_)
);

NAND2_X1 _06637_ (
  .A1(_01564_),
  .A2(din_55[7]),
  .ZN(_01571_)
);

NAND2_X1 _06638_ (
  .A1(_01570_),
  .A2(_01571_),
  .ZN(_01572_)
);

NAND2_X1 _06639_ (
  .A1(_01572_),
  .A2(_01567_),
  .ZN(_01573_)
);

NAND2_X1 _06640_ (
  .A1(_01525_),
  .A2(\sresult[12][7] ),
  .ZN(_01574_)
);

NAND2_X1 _06641_ (
  .A1(_01573_),
  .A2(_01574_),
  .ZN(_00151_)
);

BUF_X4 _06642_ (
  .A(_01519_),
  .Z(_01575_)
);

NAND2_X1 _06643_ (
  .A1(_01575_),
  .A2(\sresult[11][8] ),
  .ZN(_01576_)
);

NAND2_X1 _06644_ (
  .A1(_01564_),
  .A2(din_55[8]),
  .ZN(_01577_)
);

NAND2_X1 _06645_ (
  .A1(_01576_),
  .A2(_01577_),
  .ZN(_01578_)
);

NAND2_X1 _06646_ (
  .A1(_01578_),
  .A2(_01567_),
  .ZN(_01579_)
);

BUF_X8 _06647_ (
  .A(_00810_),
  .Z(_01580_)
);

BUF_X1 _06648_ (
  .A(_01580_),
  .Z(_01581_)
);

NAND2_X1 _06649_ (
  .A1(_01581_),
  .A2(\sresult[12][8] ),
  .ZN(_01582_)
);

NAND2_X1 _06650_ (
  .A1(_01579_),
  .A2(_01582_),
  .ZN(_00152_)
);

NAND2_X1 _06651_ (
  .A1(_01575_),
  .A2(\sresult[11][9] ),
  .ZN(_01583_)
);

NAND2_X1 _06652_ (
  .A1(_01564_),
  .A2(din_55[9]),
  .ZN(_01584_)
);

NAND2_X1 _06653_ (
  .A1(_01583_),
  .A2(_01584_),
  .ZN(_01585_)
);

NAND2_X1 _06654_ (
  .A1(_01585_),
  .A2(_01567_),
  .ZN(_01586_)
);

NAND2_X1 _06655_ (
  .A1(_01581_),
  .A2(\sresult[12][9] ),
  .ZN(_01587_)
);

NAND2_X1 _06656_ (
  .A1(_01586_),
  .A2(_01587_),
  .ZN(_00153_)
);

NAND2_X1 _06657_ (
  .A1(_01575_),
  .A2(\sresult[11][10] ),
  .ZN(_01588_)
);

NAND2_X1 _06658_ (
  .A1(_01564_),
  .A2(din_55[10]),
  .ZN(_01589_)
);

NAND2_X1 _06659_ (
  .A1(_01588_),
  .A2(_01589_),
  .ZN(_01590_)
);

NAND2_X1 _06660_ (
  .A1(_01590_),
  .A2(_01567_),
  .ZN(_01591_)
);

NAND2_X1 _06661_ (
  .A1(_01581_),
  .A2(\sresult[12][10] ),
  .ZN(_01592_)
);

NAND2_X1 _06662_ (
  .A1(_01591_),
  .A2(_01592_),
  .ZN(_00154_)
);

NAND2_X1 _06663_ (
  .A1(_01575_),
  .A2(\sresult[11][11] ),
  .ZN(_01593_)
);

NAND2_X1 _06664_ (
  .A1(_01564_),
  .A2(din_55[11]),
  .ZN(_01594_)
);

NAND2_X1 _06665_ (
  .A1(_01593_),
  .A2(_01594_),
  .ZN(_01595_)
);

NAND2_X1 _06666_ (
  .A1(_01595_),
  .A2(_01567_),
  .ZN(_01596_)
);

NAND2_X1 _06667_ (
  .A1(_01581_),
  .A2(\sresult[12][11] ),
  .ZN(_01597_)
);

NAND2_X1 _06668_ (
  .A1(_01596_),
  .A2(_01597_),
  .ZN(_00155_)
);

NAND2_X1 _06669_ (
  .A1(_01575_),
  .A2(\sresult[12][0] ),
  .ZN(_01598_)
);

NAND2_X1 _06670_ (
  .A1(_01564_),
  .A2(din_64[0]),
  .ZN(_01599_)
);

NAND2_X1 _06671_ (
  .A1(_01598_),
  .A2(_01599_),
  .ZN(_01600_)
);

NAND2_X1 _06672_ (
  .A1(_01600_),
  .A2(_01567_),
  .ZN(_01601_)
);

NAND2_X1 _06673_ (
  .A1(_01581_),
  .A2(\sresult[13][0] ),
  .ZN(_01602_)
);

NAND2_X1 _06674_ (
  .A1(_01601_),
  .A2(_01602_),
  .ZN(_00156_)
);

NAND2_X1 _06675_ (
  .A1(_01575_),
  .A2(\sresult[12][1] ),
  .ZN(_01603_)
);

NAND2_X1 _06676_ (
  .A1(_01564_),
  .A2(din_64[1]),
  .ZN(_01604_)
);

NAND2_X1 _06677_ (
  .A1(_01603_),
  .A2(_01604_),
  .ZN(_01605_)
);

NAND2_X1 _06678_ (
  .A1(_01605_),
  .A2(_01567_),
  .ZN(_01606_)
);

NAND2_X1 _06679_ (
  .A1(_01581_),
  .A2(\sresult[13][1] ),
  .ZN(_01607_)
);

NAND2_X1 _06680_ (
  .A1(_01606_),
  .A2(_01607_),
  .ZN(_00157_)
);

NAND2_X1 _06681_ (
  .A1(_01575_),
  .A2(\sresult[12][2] ),
  .ZN(_01608_)
);

NAND2_X1 _06682_ (
  .A1(_01564_),
  .A2(din_64[2]),
  .ZN(_01609_)
);

NAND2_X1 _06683_ (
  .A1(_01608_),
  .A2(_01609_),
  .ZN(_01610_)
);

NAND2_X1 _06684_ (
  .A1(_01610_),
  .A2(_01567_),
  .ZN(_01611_)
);

NAND2_X1 _06685_ (
  .A1(_01581_),
  .A2(\sresult[13][2] ),
  .ZN(_01612_)
);

NAND2_X1 _06686_ (
  .A1(_01611_),
  .A2(_01612_),
  .ZN(_00158_)
);

NAND2_X1 _06687_ (
  .A1(_01575_),
  .A2(\sresult[12][3] ),
  .ZN(_01613_)
);

NAND2_X1 _06688_ (
  .A1(_01564_),
  .A2(din_64[3]),
  .ZN(_01614_)
);

NAND2_X1 _06689_ (
  .A1(_01613_),
  .A2(_01614_),
  .ZN(_01615_)
);

NAND2_X1 _06690_ (
  .A1(_01615_),
  .A2(_01567_),
  .ZN(_01616_)
);

NAND2_X1 _06691_ (
  .A1(_01581_),
  .A2(\sresult[13][3] ),
  .ZN(_01617_)
);

NAND2_X1 _06692_ (
  .A1(_01616_),
  .A2(_01617_),
  .ZN(_00159_)
);

NAND2_X1 _06693_ (
  .A1(_01575_),
  .A2(\sresult[12][4] ),
  .ZN(_01618_)
);

BUF_X4 _06694_ (
  .A(_01563_),
  .Z(_01619_)
);

NAND2_X1 _06695_ (
  .A1(_01619_),
  .A2(din_64[4]),
  .ZN(_01620_)
);

NAND2_X1 _06696_ (
  .A1(_01618_),
  .A2(_01620_),
  .ZN(_01621_)
);

BUF_X2 _06697_ (
  .A(_01456_),
  .Z(_01622_)
);

NAND2_X1 _06698_ (
  .A1(_01621_),
  .A2(_01622_),
  .ZN(_01623_)
);

NAND2_X1 _06699_ (
  .A1(_01581_),
  .A2(\sresult[13][4] ),
  .ZN(_01624_)
);

NAND2_X1 _06700_ (
  .A1(_01623_),
  .A2(_01624_),
  .ZN(_00160_)
);

NAND2_X1 _06701_ (
  .A1(_01575_),
  .A2(\sresult[12][5] ),
  .ZN(_01625_)
);

NAND2_X1 _06702_ (
  .A1(_01619_),
  .A2(din_64[5]),
  .ZN(_01626_)
);

NAND2_X1 _06703_ (
  .A1(_01625_),
  .A2(_01626_),
  .ZN(_01627_)
);

NAND2_X1 _06704_ (
  .A1(_01627_),
  .A2(_01622_),
  .ZN(_01628_)
);

NAND2_X1 _06705_ (
  .A1(_01581_),
  .A2(\sresult[13][5] ),
  .ZN(_01629_)
);

NAND2_X1 _06706_ (
  .A1(_01628_),
  .A2(_01629_),
  .ZN(_00161_)
);

BUF_X4 _06707_ (
  .A(_01519_),
  .Z(_01630_)
);

NAND2_X1 _06708_ (
  .A1(_01630_),
  .A2(\sresult[12][6] ),
  .ZN(_01631_)
);

NAND2_X1 _06709_ (
  .A1(_01619_),
  .A2(din_64[6]),
  .ZN(_01632_)
);

NAND2_X1 _06710_ (
  .A1(_01631_),
  .A2(_01632_),
  .ZN(_01633_)
);

NAND2_X1 _06711_ (
  .A1(_01633_),
  .A2(_01622_),
  .ZN(_01634_)
);

BUF_X1 _06712_ (
  .A(_01580_),
  .Z(_01635_)
);

NAND2_X1 _06713_ (
  .A1(_01635_),
  .A2(\sresult[13][6] ),
  .ZN(_01636_)
);

NAND2_X1 _06714_ (
  .A1(_01634_),
  .A2(_01636_),
  .ZN(_00162_)
);

NAND2_X1 _06715_ (
  .A1(_01630_),
  .A2(\sresult[12][7] ),
  .ZN(_01637_)
);

NAND2_X1 _06716_ (
  .A1(_01619_),
  .A2(din_64[7]),
  .ZN(_01638_)
);

NAND2_X1 _06717_ (
  .A1(_01637_),
  .A2(_01638_),
  .ZN(_01639_)
);

NAND2_X1 _06718_ (
  .A1(_01639_),
  .A2(_01622_),
  .ZN(_01640_)
);

NAND2_X1 _06719_ (
  .A1(_01635_),
  .A2(\sresult[13][7] ),
  .ZN(_01641_)
);

NAND2_X1 _06720_ (
  .A1(_01640_),
  .A2(_01641_),
  .ZN(_00163_)
);

NAND2_X1 _06721_ (
  .A1(_01630_),
  .A2(\sresult[12][8] ),
  .ZN(_01642_)
);

NAND2_X1 _06722_ (
  .A1(_01619_),
  .A2(din_64[8]),
  .ZN(_01643_)
);

NAND2_X1 _06723_ (
  .A1(_01642_),
  .A2(_01643_),
  .ZN(_01644_)
);

NAND2_X1 _06724_ (
  .A1(_01644_),
  .A2(_01622_),
  .ZN(_01645_)
);

NAND2_X1 _06725_ (
  .A1(_01635_),
  .A2(\sresult[13][8] ),
  .ZN(_01646_)
);

NAND2_X1 _06726_ (
  .A1(_01645_),
  .A2(_01646_),
  .ZN(_00164_)
);

NAND2_X1 _06727_ (
  .A1(_01630_),
  .A2(\sresult[12][9] ),
  .ZN(_01647_)
);

NAND2_X1 _06728_ (
  .A1(_01619_),
  .A2(din_64[9]),
  .ZN(_01648_)
);

NAND2_X1 _06729_ (
  .A1(_01647_),
  .A2(_01648_),
  .ZN(_01649_)
);

NAND2_X1 _06730_ (
  .A1(_01649_),
  .A2(_01622_),
  .ZN(_01650_)
);

NAND2_X1 _06731_ (
  .A1(_01635_),
  .A2(\sresult[13][9] ),
  .ZN(_01651_)
);

NAND2_X1 _06732_ (
  .A1(_01650_),
  .A2(_01651_),
  .ZN(_00165_)
);

NAND2_X1 _06733_ (
  .A1(_01630_),
  .A2(\sresult[12][10] ),
  .ZN(_01652_)
);

NAND2_X1 _06734_ (
  .A1(_01619_),
  .A2(din_64[10]),
  .ZN(_01653_)
);

NAND2_X1 _06735_ (
  .A1(_01652_),
  .A2(_01653_),
  .ZN(_01654_)
);

NAND2_X1 _06736_ (
  .A1(_01654_),
  .A2(_01622_),
  .ZN(_01655_)
);

NAND2_X1 _06737_ (
  .A1(_01635_),
  .A2(\sresult[13][10] ),
  .ZN(_01656_)
);

NAND2_X1 _06738_ (
  .A1(_01655_),
  .A2(_01656_),
  .ZN(_00166_)
);

NAND2_X1 _06739_ (
  .A1(_01630_),
  .A2(\sresult[12][11] ),
  .ZN(_01657_)
);

NAND2_X1 _06740_ (
  .A1(_01619_),
  .A2(din_64[11]),
  .ZN(_01658_)
);

NAND2_X1 _06741_ (
  .A1(_01657_),
  .A2(_01658_),
  .ZN(_01659_)
);

NAND2_X1 _06742_ (
  .A1(_01659_),
  .A2(_01622_),
  .ZN(_01660_)
);

NAND2_X1 _06743_ (
  .A1(_01635_),
  .A2(\sresult[13][11] ),
  .ZN(_01661_)
);

NAND2_X1 _06744_ (
  .A1(_01660_),
  .A2(_01661_),
  .ZN(_00167_)
);

NAND2_X1 _06745_ (
  .A1(_01630_),
  .A2(\sresult[13][0] ),
  .ZN(_01662_)
);

NAND2_X1 _06746_ (
  .A1(_01619_),
  .A2(din_73[0]),
  .ZN(_01663_)
);

NAND2_X1 _06747_ (
  .A1(_01662_),
  .A2(_01663_),
  .ZN(_01664_)
);

NAND2_X1 _06748_ (
  .A1(_01664_),
  .A2(_01622_),
  .ZN(_01665_)
);

NAND2_X1 _06749_ (
  .A1(_01635_),
  .A2(\sresult[14][0] ),
  .ZN(_01666_)
);

NAND2_X1 _06750_ (
  .A1(_01665_),
  .A2(_01666_),
  .ZN(_00168_)
);

NAND2_X1 _06751_ (
  .A1(_01630_),
  .A2(\sresult[13][1] ),
  .ZN(_01667_)
);

NAND2_X1 _06752_ (
  .A1(_01619_),
  .A2(din_73[1]),
  .ZN(_01668_)
);

NAND2_X1 _06753_ (
  .A1(_01667_),
  .A2(_01668_),
  .ZN(_01669_)
);

NAND2_X1 _06754_ (
  .A1(_01669_),
  .A2(_01622_),
  .ZN(_01670_)
);

NAND2_X1 _06755_ (
  .A1(_01635_),
  .A2(\sresult[14][1] ),
  .ZN(_01671_)
);

NAND2_X1 _06756_ (
  .A1(_01670_),
  .A2(_01671_),
  .ZN(_00169_)
);

NAND2_X1 _06757_ (
  .A1(_01630_),
  .A2(\sresult[13][2] ),
  .ZN(_01672_)
);

BUF_X4 _06758_ (
  .A(_01563_),
  .Z(_01673_)
);

NAND2_X1 _06759_ (
  .A1(_01673_),
  .A2(din_73[2]),
  .ZN(_01674_)
);

NAND2_X1 _06760_ (
  .A1(_01672_),
  .A2(_01674_),
  .ZN(_01675_)
);

BUF_X2 _06761_ (
  .A(_01456_),
  .Z(_01676_)
);

NAND2_X1 _06762_ (
  .A1(_01675_),
  .A2(_01676_),
  .ZN(_01677_)
);

NAND2_X1 _06763_ (
  .A1(_01635_),
  .A2(\sresult[14][2] ),
  .ZN(_01678_)
);

NAND2_X1 _06764_ (
  .A1(_01677_),
  .A2(_01678_),
  .ZN(_00170_)
);

NAND2_X1 _06765_ (
  .A1(_01630_),
  .A2(\sresult[13][3] ),
  .ZN(_01679_)
);

NAND2_X1 _06766_ (
  .A1(_01673_),
  .A2(din_73[3]),
  .ZN(_01680_)
);

NAND2_X1 _06767_ (
  .A1(_01679_),
  .A2(_01680_),
  .ZN(_01681_)
);

NAND2_X1 _06768_ (
  .A1(_01681_),
  .A2(_01676_),
  .ZN(_01682_)
);

NAND2_X1 _06769_ (
  .A1(_01635_),
  .A2(\sresult[14][3] ),
  .ZN(_01683_)
);

NAND2_X1 _06770_ (
  .A1(_01682_),
  .A2(_01683_),
  .ZN(_00171_)
);

BUF_X4 _06771_ (
  .A(_01519_),
  .Z(_01684_)
);

NAND2_X1 _06772_ (
  .A1(_01684_),
  .A2(\sresult[13][4] ),
  .ZN(_01685_)
);

NAND2_X1 _06773_ (
  .A1(_01673_),
  .A2(din_73[4]),
  .ZN(_01686_)
);

NAND2_X1 _06774_ (
  .A1(_01685_),
  .A2(_01686_),
  .ZN(_01687_)
);

NAND2_X1 _06775_ (
  .A1(_01687_),
  .A2(_01676_),
  .ZN(_01688_)
);

BUF_X1 _06776_ (
  .A(_01580_),
  .Z(_01689_)
);

NAND2_X1 _06777_ (
  .A1(_01689_),
  .A2(\sresult[14][4] ),
  .ZN(_01690_)
);

NAND2_X1 _06778_ (
  .A1(_01688_),
  .A2(_01690_),
  .ZN(_00172_)
);

NAND2_X1 _06779_ (
  .A1(_01684_),
  .A2(\sresult[13][5] ),
  .ZN(_01691_)
);

NAND2_X1 _06780_ (
  .A1(_01673_),
  .A2(din_73[5]),
  .ZN(_01692_)
);

NAND2_X1 _06781_ (
  .A1(_01691_),
  .A2(_01692_),
  .ZN(_01693_)
);

NAND2_X1 _06782_ (
  .A1(_01693_),
  .A2(_01676_),
  .ZN(_01694_)
);

NAND2_X1 _06783_ (
  .A1(_01689_),
  .A2(\sresult[14][5] ),
  .ZN(_01695_)
);

NAND2_X1 _06784_ (
  .A1(_01694_),
  .A2(_01695_),
  .ZN(_00173_)
);

NAND2_X1 _06785_ (
  .A1(_01684_),
  .A2(\sresult[13][6] ),
  .ZN(_01696_)
);

NAND2_X1 _06786_ (
  .A1(_01673_),
  .A2(din_73[6]),
  .ZN(_01697_)
);

NAND2_X1 _06787_ (
  .A1(_01696_),
  .A2(_01697_),
  .ZN(_01698_)
);

NAND2_X1 _06788_ (
  .A1(_01698_),
  .A2(_01676_),
  .ZN(_01699_)
);

NAND2_X1 _06789_ (
  .A1(_01689_),
  .A2(\sresult[14][6] ),
  .ZN(_01700_)
);

NAND2_X1 _06790_ (
  .A1(_01699_),
  .A2(_01700_),
  .ZN(_00174_)
);

NAND2_X1 _06791_ (
  .A1(_01684_),
  .A2(\sresult[13][7] ),
  .ZN(_01701_)
);

NAND2_X1 _06792_ (
  .A1(_01673_),
  .A2(din_73[7]),
  .ZN(_01702_)
);

NAND2_X1 _06793_ (
  .A1(_01701_),
  .A2(_01702_),
  .ZN(_01703_)
);

NAND2_X1 _06794_ (
  .A1(_01703_),
  .A2(_01676_),
  .ZN(_01704_)
);

NAND2_X1 _06795_ (
  .A1(_01689_),
  .A2(\sresult[14][7] ),
  .ZN(_01705_)
);

NAND2_X1 _06796_ (
  .A1(_01704_),
  .A2(_01705_),
  .ZN(_00175_)
);

NAND2_X1 _06797_ (
  .A1(_01684_),
  .A2(\sresult[13][8] ),
  .ZN(_01706_)
);

NAND2_X1 _06798_ (
  .A1(_01673_),
  .A2(din_73[8]),
  .ZN(_01707_)
);

NAND2_X1 _06799_ (
  .A1(_01706_),
  .A2(_01707_),
  .ZN(_01708_)
);

NAND2_X1 _06800_ (
  .A1(_01708_),
  .A2(_01676_),
  .ZN(_01709_)
);

NAND2_X1 _06801_ (
  .A1(_01689_),
  .A2(\sresult[14][8] ),
  .ZN(_01710_)
);

NAND2_X1 _06802_ (
  .A1(_01709_),
  .A2(_01710_),
  .ZN(_00176_)
);

NAND2_X1 _06803_ (
  .A1(_01684_),
  .A2(\sresult[13][9] ),
  .ZN(_01711_)
);

NAND2_X1 _06804_ (
  .A1(_01673_),
  .A2(din_73[9]),
  .ZN(_01712_)
);

NAND2_X1 _06805_ (
  .A1(_01711_),
  .A2(_01712_),
  .ZN(_01713_)
);

NAND2_X1 _06806_ (
  .A1(_01713_),
  .A2(_01676_),
  .ZN(_01714_)
);

NAND2_X1 _06807_ (
  .A1(_01689_),
  .A2(\sresult[14][9] ),
  .ZN(_01715_)
);

NAND2_X1 _06808_ (
  .A1(_01714_),
  .A2(_01715_),
  .ZN(_00177_)
);

NAND2_X1 _06809_ (
  .A1(_01684_),
  .A2(\sresult[13][10] ),
  .ZN(_01716_)
);

NAND2_X1 _06810_ (
  .A1(_01673_),
  .A2(din_73[10]),
  .ZN(_01717_)
);

NAND2_X1 _06811_ (
  .A1(_01716_),
  .A2(_01717_),
  .ZN(_01718_)
);

NAND2_X1 _06812_ (
  .A1(_01718_),
  .A2(_01676_),
  .ZN(_01719_)
);

NAND2_X1 _06813_ (
  .A1(_01689_),
  .A2(\sresult[14][10] ),
  .ZN(_01720_)
);

NAND2_X1 _06814_ (
  .A1(_01719_),
  .A2(_01720_),
  .ZN(_00178_)
);

NAND2_X1 _06815_ (
  .A1(_01684_),
  .A2(\sresult[13][11] ),
  .ZN(_01721_)
);

NAND2_X1 _06816_ (
  .A1(_01673_),
  .A2(din_73[11]),
  .ZN(_01722_)
);

NAND2_X1 _06817_ (
  .A1(_01721_),
  .A2(_01722_),
  .ZN(_01723_)
);

NAND2_X1 _06818_ (
  .A1(_01723_),
  .A2(_01676_),
  .ZN(_01724_)
);

NAND2_X1 _06819_ (
  .A1(_01689_),
  .A2(\sresult[14][11] ),
  .ZN(_01725_)
);

NAND2_X1 _06820_ (
  .A1(_01724_),
  .A2(_01725_),
  .ZN(_00179_)
);

NAND2_X1 _06821_ (
  .A1(_01684_),
  .A2(\sresult[14][0] ),
  .ZN(_01726_)
);

BUF_X4 _06822_ (
  .A(_01563_),
  .Z(_01727_)
);

NAND2_X1 _06823_ (
  .A1(_01727_),
  .A2(din_72[0]),
  .ZN(_01728_)
);

NAND2_X1 _06824_ (
  .A1(_01726_),
  .A2(_01728_),
  .ZN(_01729_)
);

BUF_X2 _06825_ (
  .A(_01456_),
  .Z(_01730_)
);

NAND2_X1 _06826_ (
  .A1(_01729_),
  .A2(_01730_),
  .ZN(_01731_)
);

NAND2_X1 _06827_ (
  .A1(_01689_),
  .A2(\sresult[15][0] ),
  .ZN(_01732_)
);

NAND2_X1 _06828_ (
  .A1(_01731_),
  .A2(_01732_),
  .ZN(_00180_)
);

NAND2_X1 _06829_ (
  .A1(_01684_),
  .A2(\sresult[14][1] ),
  .ZN(_01733_)
);

NAND2_X1 _06830_ (
  .A1(_01727_),
  .A2(din_72[1]),
  .ZN(_01734_)
);

NAND2_X1 _06831_ (
  .A1(_01733_),
  .A2(_01734_),
  .ZN(_01735_)
);

NAND2_X1 _06832_ (
  .A1(_01735_),
  .A2(_01730_),
  .ZN(_01736_)
);

NAND2_X1 _06833_ (
  .A1(_01689_),
  .A2(\sresult[15][1] ),
  .ZN(_01737_)
);

NAND2_X1 _06834_ (
  .A1(_01736_),
  .A2(_01737_),
  .ZN(_00181_)
);

BUF_X4 _06835_ (
  .A(_01519_),
  .Z(_01738_)
);

NAND2_X1 _06836_ (
  .A1(_01738_),
  .A2(\sresult[14][2] ),
  .ZN(_01739_)
);

NAND2_X1 _06837_ (
  .A1(_01727_),
  .A2(din_72[2]),
  .ZN(_01740_)
);

NAND2_X1 _06838_ (
  .A1(_01739_),
  .A2(_01740_),
  .ZN(_01741_)
);

NAND2_X1 _06839_ (
  .A1(_01741_),
  .A2(_01730_),
  .ZN(_01742_)
);

BUF_X1 _06840_ (
  .A(_01580_),
  .Z(_01743_)
);

NAND2_X1 _06841_ (
  .A1(_01743_),
  .A2(\sresult[15][2] ),
  .ZN(_01744_)
);

NAND2_X1 _06842_ (
  .A1(_01742_),
  .A2(_01744_),
  .ZN(_00182_)
);

NAND2_X1 _06843_ (
  .A1(_01738_),
  .A2(\sresult[14][3] ),
  .ZN(_01745_)
);

NAND2_X1 _06844_ (
  .A1(_01727_),
  .A2(din_72[3]),
  .ZN(_01746_)
);

NAND2_X1 _06845_ (
  .A1(_01745_),
  .A2(_01746_),
  .ZN(_01747_)
);

NAND2_X1 _06846_ (
  .A1(_01747_),
  .A2(_01730_),
  .ZN(_01748_)
);

NAND2_X1 _06847_ (
  .A1(_01743_),
  .A2(\sresult[15][3] ),
  .ZN(_01749_)
);

NAND2_X1 _06848_ (
  .A1(_01748_),
  .A2(_01749_),
  .ZN(_00183_)
);

NAND2_X1 _06849_ (
  .A1(_01738_),
  .A2(\sresult[14][4] ),
  .ZN(_01750_)
);

NAND2_X1 _06850_ (
  .A1(_01727_),
  .A2(din_72[4]),
  .ZN(_01751_)
);

NAND2_X1 _06851_ (
  .A1(_01750_),
  .A2(_01751_),
  .ZN(_01752_)
);

NAND2_X1 _06852_ (
  .A1(_01752_),
  .A2(_01730_),
  .ZN(_01753_)
);

NAND2_X1 _06853_ (
  .A1(_01743_),
  .A2(\sresult[15][4] ),
  .ZN(_01754_)
);

NAND2_X1 _06854_ (
  .A1(_01753_),
  .A2(_01754_),
  .ZN(_00184_)
);

NAND2_X1 _06855_ (
  .A1(_01738_),
  .A2(\sresult[14][5] ),
  .ZN(_01755_)
);

NAND2_X1 _06856_ (
  .A1(_01727_),
  .A2(din_72[5]),
  .ZN(_01756_)
);

NAND2_X1 _06857_ (
  .A1(_01755_),
  .A2(_01756_),
  .ZN(_01757_)
);

NAND2_X1 _06858_ (
  .A1(_01757_),
  .A2(_01730_),
  .ZN(_01758_)
);

NAND2_X1 _06859_ (
  .A1(_01743_),
  .A2(\sresult[15][5] ),
  .ZN(_01759_)
);

NAND2_X1 _06860_ (
  .A1(_01758_),
  .A2(_01759_),
  .ZN(_00185_)
);

NAND2_X1 _06861_ (
  .A1(_01738_),
  .A2(\sresult[14][6] ),
  .ZN(_01760_)
);

NAND2_X1 _06862_ (
  .A1(_01727_),
  .A2(din_72[6]),
  .ZN(_01761_)
);

NAND2_X1 _06863_ (
  .A1(_01760_),
  .A2(_01761_),
  .ZN(_01762_)
);

NAND2_X1 _06864_ (
  .A1(_01762_),
  .A2(_01730_),
  .ZN(_01763_)
);

NAND2_X1 _06865_ (
  .A1(_01743_),
  .A2(\sresult[15][6] ),
  .ZN(_01764_)
);

NAND2_X1 _06866_ (
  .A1(_01763_),
  .A2(_01764_),
  .ZN(_00186_)
);

NAND2_X1 _06867_ (
  .A1(_01738_),
  .A2(\sresult[14][7] ),
  .ZN(_01765_)
);

NAND2_X1 _06868_ (
  .A1(_01727_),
  .A2(din_72[7]),
  .ZN(_01766_)
);

NAND2_X1 _06869_ (
  .A1(_01765_),
  .A2(_01766_),
  .ZN(_01767_)
);

NAND2_X1 _06870_ (
  .A1(_01767_),
  .A2(_01730_),
  .ZN(_01768_)
);

NAND2_X1 _06871_ (
  .A1(_01743_),
  .A2(\sresult[15][7] ),
  .ZN(_01769_)
);

NAND2_X1 _06872_ (
  .A1(_01768_),
  .A2(_01769_),
  .ZN(_00187_)
);

NAND2_X1 _06873_ (
  .A1(_01738_),
  .A2(\sresult[14][8] ),
  .ZN(_01770_)
);

NAND2_X1 _06874_ (
  .A1(_01727_),
  .A2(din_72[8]),
  .ZN(_01771_)
);

NAND2_X1 _06875_ (
  .A1(_01770_),
  .A2(_01771_),
  .ZN(_01772_)
);

NAND2_X1 _06876_ (
  .A1(_01772_),
  .A2(_01730_),
  .ZN(_01773_)
);

NAND2_X1 _06877_ (
  .A1(_01743_),
  .A2(\sresult[15][8] ),
  .ZN(_01774_)
);

NAND2_X1 _06878_ (
  .A1(_01773_),
  .A2(_01774_),
  .ZN(_00188_)
);

NAND2_X1 _06879_ (
  .A1(_01738_),
  .A2(\sresult[14][9] ),
  .ZN(_01775_)
);

NAND2_X1 _06880_ (
  .A1(_01727_),
  .A2(din_72[9]),
  .ZN(_01776_)
);

NAND2_X1 _06881_ (
  .A1(_01775_),
  .A2(_01776_),
  .ZN(_01777_)
);

NAND2_X1 _06882_ (
  .A1(_01777_),
  .A2(_01730_),
  .ZN(_01778_)
);

NAND2_X1 _06883_ (
  .A1(_01743_),
  .A2(\sresult[15][9] ),
  .ZN(_01779_)
);

NAND2_X1 _06884_ (
  .A1(_01778_),
  .A2(_01779_),
  .ZN(_00189_)
);

NAND2_X1 _06885_ (
  .A1(_01738_),
  .A2(\sresult[14][10] ),
  .ZN(_01780_)
);

BUF_X4 _06886_ (
  .A(_01563_),
  .Z(_01781_)
);

NAND2_X1 _06887_ (
  .A1(_01781_),
  .A2(din_72[10]),
  .ZN(_01782_)
);

NAND2_X1 _06888_ (
  .A1(_01780_),
  .A2(_01782_),
  .ZN(_01783_)
);

BUF_X2 _06889_ (
  .A(_01456_),
  .Z(_01784_)
);

NAND2_X1 _06890_ (
  .A1(_01783_),
  .A2(_01784_),
  .ZN(_01785_)
);

NAND2_X1 _06891_ (
  .A1(_01743_),
  .A2(\sresult[15][10] ),
  .ZN(_01786_)
);

NAND2_X1 _06892_ (
  .A1(_01785_),
  .A2(_01786_),
  .ZN(_00190_)
);

NAND2_X1 _06893_ (
  .A1(_01738_),
  .A2(\sresult[14][11] ),
  .ZN(_01787_)
);

NAND2_X1 _06894_ (
  .A1(_01781_),
  .A2(din_72[11]),
  .ZN(_01788_)
);

NAND2_X1 _06895_ (
  .A1(_01787_),
  .A2(_01788_),
  .ZN(_01789_)
);

NAND2_X1 _06896_ (
  .A1(_01789_),
  .A2(_01784_),
  .ZN(_01790_)
);

NAND2_X1 _06897_ (
  .A1(_01743_),
  .A2(\sresult[15][11] ),
  .ZN(_01791_)
);

NAND2_X1 _06898_ (
  .A1(_01790_),
  .A2(_01791_),
  .ZN(_00191_)
);

BUF_X4 _06899_ (
  .A(_01519_),
  .Z(_01792_)
);

NAND2_X1 _06900_ (
  .A1(_01792_),
  .A2(\sresult[15][0] ),
  .ZN(_01793_)
);

NAND2_X1 _06901_ (
  .A1(_01781_),
  .A2(din_63[0]),
  .ZN(_01794_)
);

NAND2_X1 _06902_ (
  .A1(_01793_),
  .A2(_01794_),
  .ZN(_01795_)
);

NAND2_X1 _06903_ (
  .A1(_01795_),
  .A2(_01784_),
  .ZN(_01796_)
);

BUF_X1 _06904_ (
  .A(_01580_),
  .Z(_01797_)
);

NAND2_X1 _06905_ (
  .A1(_01797_),
  .A2(\sresult[16][0] ),
  .ZN(_01798_)
);

NAND2_X1 _06906_ (
  .A1(_01796_),
  .A2(_01798_),
  .ZN(_00192_)
);

NAND2_X1 _06907_ (
  .A1(_01792_),
  .A2(\sresult[15][1] ),
  .ZN(_01799_)
);

NAND2_X1 _06908_ (
  .A1(_01781_),
  .A2(din_63[1]),
  .ZN(_01800_)
);

NAND2_X1 _06909_ (
  .A1(_01799_),
  .A2(_01800_),
  .ZN(_01801_)
);

NAND2_X1 _06910_ (
  .A1(_01801_),
  .A2(_01784_),
  .ZN(_01802_)
);

NAND2_X1 _06911_ (
  .A1(_01797_),
  .A2(\sresult[16][1] ),
  .ZN(_01803_)
);

NAND2_X1 _06912_ (
  .A1(_01802_),
  .A2(_01803_),
  .ZN(_00193_)
);

NAND2_X1 _06913_ (
  .A1(_01792_),
  .A2(\sresult[15][2] ),
  .ZN(_01804_)
);

NAND2_X1 _06914_ (
  .A1(_01781_),
  .A2(din_63[2]),
  .ZN(_01805_)
);

NAND2_X1 _06915_ (
  .A1(_01804_),
  .A2(_01805_),
  .ZN(_01806_)
);

NAND2_X1 _06916_ (
  .A1(_01806_),
  .A2(_01784_),
  .ZN(_01807_)
);

NAND2_X1 _06917_ (
  .A1(_01797_),
  .A2(\sresult[16][2] ),
  .ZN(_01808_)
);

NAND2_X1 _06918_ (
  .A1(_01807_),
  .A2(_01808_),
  .ZN(_00194_)
);

NAND2_X1 _06919_ (
  .A1(_01792_),
  .A2(\sresult[15][3] ),
  .ZN(_01809_)
);

NAND2_X1 _06920_ (
  .A1(_01781_),
  .A2(din_63[3]),
  .ZN(_01810_)
);

NAND2_X1 _06921_ (
  .A1(_01809_),
  .A2(_01810_),
  .ZN(_01811_)
);

NAND2_X1 _06922_ (
  .A1(_01811_),
  .A2(_01784_),
  .ZN(_01812_)
);

NAND2_X1 _06923_ (
  .A1(_01797_),
  .A2(\sresult[16][3] ),
  .ZN(_01813_)
);

NAND2_X1 _06924_ (
  .A1(_01812_),
  .A2(_01813_),
  .ZN(_00195_)
);

NAND2_X1 _06925_ (
  .A1(_01792_),
  .A2(\sresult[15][4] ),
  .ZN(_01814_)
);

NAND2_X1 _06926_ (
  .A1(_01781_),
  .A2(din_63[4]),
  .ZN(_01815_)
);

NAND2_X1 _06927_ (
  .A1(_01814_),
  .A2(_01815_),
  .ZN(_01816_)
);

NAND2_X1 _06928_ (
  .A1(_01816_),
  .A2(_01784_),
  .ZN(_01817_)
);

NAND2_X1 _06929_ (
  .A1(_01797_),
  .A2(\sresult[16][4] ),
  .ZN(_01818_)
);

NAND2_X1 _06930_ (
  .A1(_01817_),
  .A2(_01818_),
  .ZN(_00196_)
);

NAND2_X1 _06931_ (
  .A1(_01792_),
  .A2(\sresult[15][5] ),
  .ZN(_01819_)
);

NAND2_X1 _06932_ (
  .A1(_01781_),
  .A2(din_63[5]),
  .ZN(_01820_)
);

NAND2_X1 _06933_ (
  .A1(_01819_),
  .A2(_01820_),
  .ZN(_01821_)
);

NAND2_X1 _06934_ (
  .A1(_01821_),
  .A2(_01784_),
  .ZN(_01822_)
);

NAND2_X1 _06935_ (
  .A1(_01797_),
  .A2(\sresult[16][5] ),
  .ZN(_01823_)
);

NAND2_X1 _06936_ (
  .A1(_01822_),
  .A2(_01823_),
  .ZN(_00197_)
);

NAND2_X1 _06937_ (
  .A1(_01792_),
  .A2(\sresult[15][6] ),
  .ZN(_01824_)
);

NAND2_X1 _06938_ (
  .A1(_01781_),
  .A2(din_63[6]),
  .ZN(_01825_)
);

NAND2_X1 _06939_ (
  .A1(_01824_),
  .A2(_01825_),
  .ZN(_01826_)
);

NAND2_X1 _06940_ (
  .A1(_01826_),
  .A2(_01784_),
  .ZN(_01827_)
);

NAND2_X1 _06941_ (
  .A1(_01797_),
  .A2(\sresult[16][6] ),
  .ZN(_01828_)
);

NAND2_X1 _06942_ (
  .A1(_01827_),
  .A2(_01828_),
  .ZN(_00198_)
);

NAND2_X1 _06943_ (
  .A1(_01792_),
  .A2(\sresult[15][7] ),
  .ZN(_01829_)
);

NAND2_X1 _06944_ (
  .A1(_01781_),
  .A2(din_63[7]),
  .ZN(_01830_)
);

NAND2_X1 _06945_ (
  .A1(_01829_),
  .A2(_01830_),
  .ZN(_01831_)
);

NAND2_X1 _06946_ (
  .A1(_01831_),
  .A2(_01784_),
  .ZN(_01832_)
);

NAND2_X1 _06947_ (
  .A1(_01797_),
  .A2(\sresult[16][7] ),
  .ZN(_01833_)
);

NAND2_X1 _06948_ (
  .A1(_01832_),
  .A2(_01833_),
  .ZN(_00199_)
);

NAND2_X1 _06949_ (
  .A1(_01792_),
  .A2(\sresult[15][8] ),
  .ZN(_01834_)
);

BUF_X4 _06950_ (
  .A(_01563_),
  .Z(_01835_)
);

NAND2_X1 _06951_ (
  .A1(_01835_),
  .A2(din_63[8]),
  .ZN(_01836_)
);

NAND2_X1 _06952_ (
  .A1(_01834_),
  .A2(_01836_),
  .ZN(_01837_)
);

BUF_X2 _06953_ (
  .A(_01456_),
  .Z(_01838_)
);

NAND2_X1 _06954_ (
  .A1(_01837_),
  .A2(_01838_),
  .ZN(_01839_)
);

NAND2_X1 _06955_ (
  .A1(_01797_),
  .A2(\sresult[16][8] ),
  .ZN(_01840_)
);

NAND2_X1 _06956_ (
  .A1(_01839_),
  .A2(_01840_),
  .ZN(_00200_)
);

NAND2_X1 _06957_ (
  .A1(_01792_),
  .A2(\sresult[15][9] ),
  .ZN(_01841_)
);

NAND2_X1 _06958_ (
  .A1(_01835_),
  .A2(din_63[9]),
  .ZN(_01842_)
);

NAND2_X1 _06959_ (
  .A1(_01841_),
  .A2(_01842_),
  .ZN(_01843_)
);

NAND2_X1 _06960_ (
  .A1(_01843_),
  .A2(_01838_),
  .ZN(_01844_)
);

NAND2_X1 _06961_ (
  .A1(_01797_),
  .A2(\sresult[16][9] ),
  .ZN(_01845_)
);

NAND2_X1 _06962_ (
  .A1(_01844_),
  .A2(_01845_),
  .ZN(_00201_)
);

BUF_X4 _06963_ (
  .A(_01519_),
  .Z(_01846_)
);

NAND2_X1 _06964_ (
  .A1(_01846_),
  .A2(\sresult[15][10] ),
  .ZN(_01847_)
);

NAND2_X1 _06965_ (
  .A1(_01835_),
  .A2(din_63[10]),
  .ZN(_01848_)
);

NAND2_X1 _06966_ (
  .A1(_01847_),
  .A2(_01848_),
  .ZN(_01849_)
);

NAND2_X1 _06967_ (
  .A1(_01849_),
  .A2(_01838_),
  .ZN(_01850_)
);

BUF_X1 _06968_ (
  .A(_01580_),
  .Z(_01851_)
);

NAND2_X1 _06969_ (
  .A1(_01851_),
  .A2(\sresult[16][10] ),
  .ZN(_01852_)
);

NAND2_X1 _06970_ (
  .A1(_01850_),
  .A2(_01852_),
  .ZN(_00202_)
);

NAND2_X1 _06971_ (
  .A1(_01846_),
  .A2(\sresult[15][11] ),
  .ZN(_01853_)
);

NAND2_X1 _06972_ (
  .A1(_01835_),
  .A2(din_63[11]),
  .ZN(_01854_)
);

NAND2_X1 _06973_ (
  .A1(_01853_),
  .A2(_01854_),
  .ZN(_01855_)
);

NAND2_X1 _06974_ (
  .A1(_01855_),
  .A2(_01838_),
  .ZN(_01856_)
);

NAND2_X1 _06975_ (
  .A1(_01851_),
  .A2(\sresult[16][11] ),
  .ZN(_01857_)
);

NAND2_X1 _06976_ (
  .A1(_01856_),
  .A2(_01857_),
  .ZN(_00203_)
);

NAND2_X1 _06977_ (
  .A1(_01846_),
  .A2(\sresult[16][0] ),
  .ZN(_01858_)
);

NAND2_X1 _06978_ (
  .A1(_01835_),
  .A2(din_54[0]),
  .ZN(_01859_)
);

NAND2_X1 _06979_ (
  .A1(_01858_),
  .A2(_01859_),
  .ZN(_01860_)
);

NAND2_X1 _06980_ (
  .A1(_01860_),
  .A2(_01838_),
  .ZN(_01861_)
);

NAND2_X1 _06981_ (
  .A1(_01851_),
  .A2(\sresult[17][0] ),
  .ZN(_01862_)
);

NAND2_X1 _06982_ (
  .A1(_01861_),
  .A2(_01862_),
  .ZN(_00204_)
);

NAND2_X1 _06983_ (
  .A1(_01846_),
  .A2(\sresult[16][1] ),
  .ZN(_01863_)
);

NAND2_X1 _06984_ (
  .A1(_01835_),
  .A2(din_54[1]),
  .ZN(_01864_)
);

NAND2_X1 _06985_ (
  .A1(_01863_),
  .A2(_01864_),
  .ZN(_01865_)
);

NAND2_X1 _06986_ (
  .A1(_01865_),
  .A2(_01838_),
  .ZN(_01866_)
);

NAND2_X1 _06987_ (
  .A1(_01851_),
  .A2(\sresult[17][1] ),
  .ZN(_01867_)
);

NAND2_X1 _06988_ (
  .A1(_01866_),
  .A2(_01867_),
  .ZN(_00205_)
);

NAND2_X1 _06989_ (
  .A1(_01846_),
  .A2(\sresult[16][2] ),
  .ZN(_01868_)
);

NAND2_X1 _06990_ (
  .A1(_01835_),
  .A2(din_54[2]),
  .ZN(_01869_)
);

NAND2_X1 _06991_ (
  .A1(_01868_),
  .A2(_01869_),
  .ZN(_01870_)
);

NAND2_X1 _06992_ (
  .A1(_01870_),
  .A2(_01838_),
  .ZN(_01871_)
);

NAND2_X1 _06993_ (
  .A1(_01851_),
  .A2(\sresult[17][2] ),
  .ZN(_01872_)
);

NAND2_X1 _06994_ (
  .A1(_01871_),
  .A2(_01872_),
  .ZN(_00206_)
);

NAND2_X1 _06995_ (
  .A1(_01846_),
  .A2(\sresult[16][3] ),
  .ZN(_01873_)
);

NAND2_X1 _06996_ (
  .A1(_01835_),
  .A2(din_54[3]),
  .ZN(_01874_)
);

NAND2_X1 _06997_ (
  .A1(_01873_),
  .A2(_01874_),
  .ZN(_01875_)
);

NAND2_X1 _06998_ (
  .A1(_01875_),
  .A2(_01838_),
  .ZN(_01876_)
);

NAND2_X1 _06999_ (
  .A1(_01851_),
  .A2(\sresult[17][3] ),
  .ZN(_01877_)
);

NAND2_X1 _07000_ (
  .A1(_01876_),
  .A2(_01877_),
  .ZN(_00207_)
);

NAND2_X1 _07001_ (
  .A1(_01846_),
  .A2(\sresult[16][4] ),
  .ZN(_01878_)
);

NAND2_X1 _07002_ (
  .A1(_01835_),
  .A2(din_54[4]),
  .ZN(_01879_)
);

NAND2_X1 _07003_ (
  .A1(_01878_),
  .A2(_01879_),
  .ZN(_01880_)
);

NAND2_X1 _07004_ (
  .A1(_01880_),
  .A2(_01838_),
  .ZN(_01881_)
);

NAND2_X1 _07005_ (
  .A1(_01851_),
  .A2(\sresult[17][4] ),
  .ZN(_01882_)
);

NAND2_X1 _07006_ (
  .A1(_01881_),
  .A2(_01882_),
  .ZN(_00208_)
);

NAND2_X1 _07007_ (
  .A1(_01846_),
  .A2(\sresult[16][5] ),
  .ZN(_01883_)
);

NAND2_X1 _07008_ (
  .A1(_01835_),
  .A2(din_54[5]),
  .ZN(_01884_)
);

NAND2_X1 _07009_ (
  .A1(_01883_),
  .A2(_01884_),
  .ZN(_01885_)
);

NAND2_X1 _07010_ (
  .A1(_01885_),
  .A2(_01838_),
  .ZN(_01886_)
);

NAND2_X1 _07011_ (
  .A1(_01851_),
  .A2(\sresult[17][5] ),
  .ZN(_01887_)
);

NAND2_X1 _07012_ (
  .A1(_01886_),
  .A2(_01887_),
  .ZN(_00209_)
);

NAND2_X1 _07013_ (
  .A1(_01846_),
  .A2(\sresult[16][6] ),
  .ZN(_01888_)
);

BUF_X4 _07014_ (
  .A(_01563_),
  .Z(_01889_)
);

NAND2_X1 _07015_ (
  .A1(_01889_),
  .A2(din_54[6]),
  .ZN(_01890_)
);

NAND2_X1 _07016_ (
  .A1(_01888_),
  .A2(_01890_),
  .ZN(_01891_)
);

BUF_X2 _07017_ (
  .A(_01456_),
  .Z(_01892_)
);

NAND2_X1 _07018_ (
  .A1(_01891_),
  .A2(_01892_),
  .ZN(_01893_)
);

NAND2_X1 _07019_ (
  .A1(_01851_),
  .A2(\sresult[17][6] ),
  .ZN(_01894_)
);

NAND2_X1 _07020_ (
  .A1(_01893_),
  .A2(_01894_),
  .ZN(_00210_)
);

NAND2_X1 _07021_ (
  .A1(_01846_),
  .A2(\sresult[16][7] ),
  .ZN(_01895_)
);

NAND2_X1 _07022_ (
  .A1(_01889_),
  .A2(din_54[7]),
  .ZN(_01896_)
);

NAND2_X1 _07023_ (
  .A1(_01895_),
  .A2(_01896_),
  .ZN(_01897_)
);

NAND2_X1 _07024_ (
  .A1(_01897_),
  .A2(_01892_),
  .ZN(_01898_)
);

NAND2_X1 _07025_ (
  .A1(_01851_),
  .A2(\sresult[17][7] ),
  .ZN(_01899_)
);

NAND2_X1 _07026_ (
  .A1(_01898_),
  .A2(_01899_),
  .ZN(_00211_)
);

BUF_X4 _07027_ (
  .A(_01519_),
  .Z(_01900_)
);

NAND2_X1 _07028_ (
  .A1(_01900_),
  .A2(\sresult[16][8] ),
  .ZN(_01901_)
);

NAND2_X1 _07029_ (
  .A1(_01889_),
  .A2(din_54[8]),
  .ZN(_01902_)
);

NAND2_X1 _07030_ (
  .A1(_01901_),
  .A2(_01902_),
  .ZN(_01903_)
);

NAND2_X1 _07031_ (
  .A1(_01903_),
  .A2(_01892_),
  .ZN(_01904_)
);

BUF_X1 _07032_ (
  .A(_01580_),
  .Z(_01905_)
);

NAND2_X1 _07033_ (
  .A1(_01905_),
  .A2(\sresult[17][8] ),
  .ZN(_01906_)
);

NAND2_X1 _07034_ (
  .A1(_01904_),
  .A2(_01906_),
  .ZN(_00212_)
);

NAND2_X1 _07035_ (
  .A1(_01900_),
  .A2(\sresult[16][9] ),
  .ZN(_01907_)
);

NAND2_X1 _07036_ (
  .A1(_01889_),
  .A2(din_54[9]),
  .ZN(_01908_)
);

NAND2_X1 _07037_ (
  .A1(_01907_),
  .A2(_01908_),
  .ZN(_01909_)
);

NAND2_X1 _07038_ (
  .A1(_01909_),
  .A2(_01892_),
  .ZN(_01910_)
);

NAND2_X1 _07039_ (
  .A1(_01905_),
  .A2(\sresult[17][9] ),
  .ZN(_01911_)
);

NAND2_X1 _07040_ (
  .A1(_01910_),
  .A2(_01911_),
  .ZN(_00213_)
);

NAND2_X1 _07041_ (
  .A1(_01900_),
  .A2(\sresult[16][10] ),
  .ZN(_01912_)
);

NAND2_X1 _07042_ (
  .A1(_01889_),
  .A2(din_54[10]),
  .ZN(_01913_)
);

NAND2_X1 _07043_ (
  .A1(_01912_),
  .A2(_01913_),
  .ZN(_01914_)
);

NAND2_X1 _07044_ (
  .A1(_01914_),
  .A2(_01892_),
  .ZN(_01915_)
);

NAND2_X1 _07045_ (
  .A1(_01905_),
  .A2(\sresult[17][10] ),
  .ZN(_01916_)
);

NAND2_X1 _07046_ (
  .A1(_01915_),
  .A2(_01916_),
  .ZN(_00214_)
);

NAND2_X1 _07047_ (
  .A1(_01900_),
  .A2(\sresult[16][11] ),
  .ZN(_01917_)
);

NAND2_X1 _07048_ (
  .A1(_01889_),
  .A2(din_54[11]),
  .ZN(_01918_)
);

NAND2_X1 _07049_ (
  .A1(_01917_),
  .A2(_01918_),
  .ZN(_01919_)
);

NAND2_X1 _07050_ (
  .A1(_01919_),
  .A2(_01892_),
  .ZN(_01920_)
);

NAND2_X1 _07051_ (
  .A1(_01905_),
  .A2(\sresult[17][11] ),
  .ZN(_01921_)
);

NAND2_X1 _07052_ (
  .A1(_01920_),
  .A2(_01921_),
  .ZN(_00215_)
);

NAND2_X1 _07053_ (
  .A1(_01900_),
  .A2(\sresult[17][0] ),
  .ZN(_01922_)
);

NAND2_X1 _07054_ (
  .A1(_01889_),
  .A2(din_45[0]),
  .ZN(_01923_)
);

NAND2_X1 _07055_ (
  .A1(_01922_),
  .A2(_01923_),
  .ZN(_01924_)
);

NAND2_X1 _07056_ (
  .A1(_01924_),
  .A2(_01892_),
  .ZN(_01925_)
);

NAND2_X1 _07057_ (
  .A1(_01905_),
  .A2(\sresult[18][0] ),
  .ZN(_01926_)
);

NAND2_X1 _07058_ (
  .A1(_01925_),
  .A2(_01926_),
  .ZN(_00216_)
);

NAND2_X1 _07059_ (
  .A1(_01900_),
  .A2(\sresult[17][1] ),
  .ZN(_01927_)
);

NAND2_X1 _07060_ (
  .A1(_01889_),
  .A2(din_45[1]),
  .ZN(_01928_)
);

NAND2_X1 _07061_ (
  .A1(_01927_),
  .A2(_01928_),
  .ZN(_01929_)
);

NAND2_X1 _07062_ (
  .A1(_01929_),
  .A2(_01892_),
  .ZN(_01930_)
);

NAND2_X1 _07063_ (
  .A1(_01905_),
  .A2(\sresult[18][1] ),
  .ZN(_01931_)
);

NAND2_X1 _07064_ (
  .A1(_01930_),
  .A2(_01931_),
  .ZN(_00217_)
);

NAND2_X1 _07065_ (
  .A1(_01900_),
  .A2(\sresult[17][2] ),
  .ZN(_01932_)
);

NAND2_X1 _07066_ (
  .A1(_01889_),
  .A2(din_45[2]),
  .ZN(_01933_)
);

NAND2_X1 _07067_ (
  .A1(_01932_),
  .A2(_01933_),
  .ZN(_01934_)
);

NAND2_X1 _07068_ (
  .A1(_01934_),
  .A2(_01892_),
  .ZN(_01935_)
);

NAND2_X1 _07069_ (
  .A1(_01905_),
  .A2(\sresult[18][2] ),
  .ZN(_01936_)
);

NAND2_X1 _07070_ (
  .A1(_01935_),
  .A2(_01936_),
  .ZN(_00218_)
);

NAND2_X1 _07071_ (
  .A1(_01900_),
  .A2(\sresult[17][3] ),
  .ZN(_01937_)
);

NAND2_X1 _07072_ (
  .A1(_01889_),
  .A2(din_45[3]),
  .ZN(_01938_)
);

NAND2_X1 _07073_ (
  .A1(_01937_),
  .A2(_01938_),
  .ZN(_01939_)
);

NAND2_X1 _07074_ (
  .A1(_01939_),
  .A2(_01892_),
  .ZN(_01940_)
);

NAND2_X1 _07075_ (
  .A1(_01905_),
  .A2(\sresult[18][3] ),
  .ZN(_01941_)
);

NAND2_X1 _07076_ (
  .A1(_01940_),
  .A2(_01941_),
  .ZN(_00219_)
);

NAND2_X1 _07077_ (
  .A1(_01900_),
  .A2(\sresult[17][4] ),
  .ZN(_01942_)
);

BUF_X4 _07078_ (
  .A(_01563_),
  .Z(_01943_)
);

NAND2_X1 _07079_ (
  .A1(_01943_),
  .A2(din_45[4]),
  .ZN(_01944_)
);

NAND2_X1 _07080_ (
  .A1(_01942_),
  .A2(_01944_),
  .ZN(_01945_)
);

BUF_X2 _07081_ (
  .A(_01456_),
  .Z(_01946_)
);

NAND2_X1 _07082_ (
  .A1(_01945_),
  .A2(_01946_),
  .ZN(_01947_)
);

NAND2_X1 _07083_ (
  .A1(_01905_),
  .A2(\sresult[18][4] ),
  .ZN(_01948_)
);

NAND2_X1 _07084_ (
  .A1(_01947_),
  .A2(_01948_),
  .ZN(_00220_)
);

NAND2_X1 _07085_ (
  .A1(_01900_),
  .A2(\sresult[17][5] ),
  .ZN(_01949_)
);

NAND2_X1 _07086_ (
  .A1(_01943_),
  .A2(din_45[5]),
  .ZN(_01950_)
);

NAND2_X1 _07087_ (
  .A1(_01949_),
  .A2(_01950_),
  .ZN(_01951_)
);

NAND2_X1 _07088_ (
  .A1(_01951_),
  .A2(_01946_),
  .ZN(_01952_)
);

NAND2_X1 _07089_ (
  .A1(_01905_),
  .A2(\sresult[18][5] ),
  .ZN(_01953_)
);

NAND2_X1 _07090_ (
  .A1(_01952_),
  .A2(_01953_),
  .ZN(_00221_)
);

BUF_X4 _07091_ (
  .A(_01519_),
  .Z(_01954_)
);

NAND2_X1 _07092_ (
  .A1(_01954_),
  .A2(\sresult[17][6] ),
  .ZN(_01955_)
);

NAND2_X1 _07093_ (
  .A1(_01943_),
  .A2(din_45[6]),
  .ZN(_01956_)
);

NAND2_X1 _07094_ (
  .A1(_01955_),
  .A2(_01956_),
  .ZN(_01957_)
);

NAND2_X1 _07095_ (
  .A1(_01957_),
  .A2(_01946_),
  .ZN(_01958_)
);

BUF_X1 _07096_ (
  .A(_01580_),
  .Z(_01959_)
);

NAND2_X1 _07097_ (
  .A1(_01959_),
  .A2(\sresult[18][6] ),
  .ZN(_01960_)
);

NAND2_X1 _07098_ (
  .A1(_01958_),
  .A2(_01960_),
  .ZN(_00222_)
);

NAND2_X1 _07099_ (
  .A1(_01954_),
  .A2(\sresult[17][7] ),
  .ZN(_01961_)
);

NAND2_X1 _07100_ (
  .A1(_01943_),
  .A2(din_45[7]),
  .ZN(_01962_)
);

NAND2_X1 _07101_ (
  .A1(_01961_),
  .A2(_01962_),
  .ZN(_01963_)
);

NAND2_X1 _07102_ (
  .A1(_01963_),
  .A2(_01946_),
  .ZN(_01964_)
);

NAND2_X1 _07103_ (
  .A1(_01959_),
  .A2(\sresult[18][7] ),
  .ZN(_01965_)
);

NAND2_X1 _07104_ (
  .A1(_01964_),
  .A2(_01965_),
  .ZN(_00223_)
);

NAND2_X1 _07105_ (
  .A1(_01954_),
  .A2(\sresult[17][8] ),
  .ZN(_01966_)
);

NAND2_X1 _07106_ (
  .A1(_01943_),
  .A2(din_45[8]),
  .ZN(_01967_)
);

NAND2_X1 _07107_ (
  .A1(_01966_),
  .A2(_01967_),
  .ZN(_01968_)
);

NAND2_X1 _07108_ (
  .A1(_01968_),
  .A2(_01946_),
  .ZN(_01969_)
);

NAND2_X1 _07109_ (
  .A1(_01959_),
  .A2(\sresult[18][8] ),
  .ZN(_01970_)
);

NAND2_X1 _07110_ (
  .A1(_01969_),
  .A2(_01970_),
  .ZN(_00224_)
);

NAND2_X1 _07111_ (
  .A1(_01954_),
  .A2(\sresult[17][9] ),
  .ZN(_01971_)
);

NAND2_X1 _07112_ (
  .A1(_01943_),
  .A2(din_45[9]),
  .ZN(_01972_)
);

NAND2_X1 _07113_ (
  .A1(_01971_),
  .A2(_01972_),
  .ZN(_01973_)
);

NAND2_X1 _07114_ (
  .A1(_01973_),
  .A2(_01946_),
  .ZN(_01974_)
);

NAND2_X1 _07115_ (
  .A1(_01959_),
  .A2(\sresult[18][9] ),
  .ZN(_01975_)
);

NAND2_X1 _07116_ (
  .A1(_01974_),
  .A2(_01975_),
  .ZN(_00225_)
);

NAND2_X1 _07117_ (
  .A1(_01954_),
  .A2(\sresult[17][10] ),
  .ZN(_01976_)
);

NAND2_X1 _07118_ (
  .A1(_01943_),
  .A2(din_45[10]),
  .ZN(_01977_)
);

NAND2_X1 _07119_ (
  .A1(_01976_),
  .A2(_01977_),
  .ZN(_01978_)
);

NAND2_X1 _07120_ (
  .A1(_01978_),
  .A2(_01946_),
  .ZN(_01979_)
);

NAND2_X1 _07121_ (
  .A1(_01959_),
  .A2(\sresult[18][10] ),
  .ZN(_01980_)
);

NAND2_X1 _07122_ (
  .A1(_01979_),
  .A2(_01980_),
  .ZN(_00226_)
);

NAND2_X1 _07123_ (
  .A1(_01954_),
  .A2(\sresult[17][11] ),
  .ZN(_01981_)
);

NAND2_X1 _07124_ (
  .A1(_01943_),
  .A2(din_45[11]),
  .ZN(_01982_)
);

NAND2_X1 _07125_ (
  .A1(_01981_),
  .A2(_01982_),
  .ZN(_01983_)
);

NAND2_X1 _07126_ (
  .A1(_01983_),
  .A2(_01946_),
  .ZN(_01984_)
);

NAND2_X1 _07127_ (
  .A1(_01959_),
  .A2(\sresult[18][11] ),
  .ZN(_01985_)
);

NAND2_X1 _07128_ (
  .A1(_01984_),
  .A2(_01985_),
  .ZN(_00227_)
);

NAND2_X1 _07129_ (
  .A1(_01954_),
  .A2(\sresult[18][0] ),
  .ZN(_01986_)
);

NAND2_X1 _07130_ (
  .A1(_01943_),
  .A2(din_36[0]),
  .ZN(_01987_)
);

NAND2_X1 _07131_ (
  .A1(_01986_),
  .A2(_01987_),
  .ZN(_01988_)
);

NAND2_X1 _07132_ (
  .A1(_01988_),
  .A2(_01946_),
  .ZN(_01989_)
);

NAND2_X1 _07133_ (
  .A1(_01959_),
  .A2(\sresult[19][0] ),
  .ZN(_01990_)
);

NAND2_X1 _07134_ (
  .A1(_01989_),
  .A2(_01990_),
  .ZN(_00228_)
);

NAND2_X1 _07135_ (
  .A1(_01954_),
  .A2(\sresult[18][1] ),
  .ZN(_01991_)
);

NAND2_X1 _07136_ (
  .A1(_01943_),
  .A2(din_36[1]),
  .ZN(_01992_)
);

NAND2_X1 _07137_ (
  .A1(_01991_),
  .A2(_01992_),
  .ZN(_01993_)
);

NAND2_X1 _07138_ (
  .A1(_01993_),
  .A2(_01946_),
  .ZN(_01994_)
);

NAND2_X1 _07139_ (
  .A1(_01959_),
  .A2(\sresult[19][1] ),
  .ZN(_01995_)
);

NAND2_X1 _07140_ (
  .A1(_01994_),
  .A2(_01995_),
  .ZN(_00229_)
);

NAND2_X1 _07141_ (
  .A1(_01954_),
  .A2(\sresult[18][2] ),
  .ZN(_01996_)
);

BUF_X4 _07142_ (
  .A(_01563_),
  .Z(_01997_)
);

NAND2_X1 _07143_ (
  .A1(_01997_),
  .A2(din_36[2]),
  .ZN(_01998_)
);

NAND2_X1 _07144_ (
  .A1(_01996_),
  .A2(_01998_),
  .ZN(_01999_)
);

BUF_X4 _07145_ (
  .A(_00911_),
  .Z(_02000_)
);

BUF_X2 _07146_ (
  .A(_02000_),
  .Z(_02001_)
);

NAND2_X1 _07147_ (
  .A1(_01999_),
  .A2(_02001_),
  .ZN(_02002_)
);

NAND2_X1 _07148_ (
  .A1(_01959_),
  .A2(\sresult[19][2] ),
  .ZN(_02003_)
);

NAND2_X1 _07149_ (
  .A1(_02002_),
  .A2(_02003_),
  .ZN(_00230_)
);

NAND2_X1 _07150_ (
  .A1(_01954_),
  .A2(\sresult[18][3] ),
  .ZN(_02004_)
);

NAND2_X1 _07151_ (
  .A1(_01997_),
  .A2(din_36[3]),
  .ZN(_02005_)
);

NAND2_X1 _07152_ (
  .A1(_02004_),
  .A2(_02005_),
  .ZN(_02006_)
);

NAND2_X1 _07153_ (
  .A1(_02006_),
  .A2(_02001_),
  .ZN(_02007_)
);

NAND2_X1 _07154_ (
  .A1(_01959_),
  .A2(\sresult[19][3] ),
  .ZN(_02008_)
);

NAND2_X1 _07155_ (
  .A1(_02007_),
  .A2(_02008_),
  .ZN(_00231_)
);

BUF_X4 _07156_ (
  .A(_01519_),
  .Z(_02009_)
);

NAND2_X1 _07157_ (
  .A1(_02009_),
  .A2(\sresult[18][4] ),
  .ZN(_02010_)
);

NAND2_X1 _07158_ (
  .A1(_01997_),
  .A2(din_36[4]),
  .ZN(_02011_)
);

NAND2_X1 _07159_ (
  .A1(_02010_),
  .A2(_02011_),
  .ZN(_02012_)
);

NAND2_X1 _07160_ (
  .A1(_02012_),
  .A2(_02001_),
  .ZN(_02013_)
);

BUF_X1 _07161_ (
  .A(_01580_),
  .Z(_02014_)
);

NAND2_X1 _07162_ (
  .A1(_02014_),
  .A2(\sresult[19][4] ),
  .ZN(_02015_)
);

NAND2_X1 _07163_ (
  .A1(_02013_),
  .A2(_02015_),
  .ZN(_00232_)
);

NAND2_X1 _07164_ (
  .A1(_02009_),
  .A2(\sresult[18][5] ),
  .ZN(_02016_)
);

NAND2_X1 _07165_ (
  .A1(_01997_),
  .A2(din_36[5]),
  .ZN(_02017_)
);

NAND2_X1 _07166_ (
  .A1(_02016_),
  .A2(_02017_),
  .ZN(_02018_)
);

NAND2_X1 _07167_ (
  .A1(_02018_),
  .A2(_02001_),
  .ZN(_02019_)
);

NAND2_X1 _07168_ (
  .A1(_02014_),
  .A2(\sresult[19][5] ),
  .ZN(_02020_)
);

NAND2_X1 _07169_ (
  .A1(_02019_),
  .A2(_02020_),
  .ZN(_00233_)
);

NAND2_X1 _07170_ (
  .A1(_02009_),
  .A2(\sresult[18][6] ),
  .ZN(_02021_)
);

NAND2_X1 _07171_ (
  .A1(_01997_),
  .A2(din_36[6]),
  .ZN(_02022_)
);

NAND2_X1 _07172_ (
  .A1(_02021_),
  .A2(_02022_),
  .ZN(_02023_)
);

NAND2_X1 _07173_ (
  .A1(_02023_),
  .A2(_02001_),
  .ZN(_02024_)
);

NAND2_X1 _07174_ (
  .A1(_02014_),
  .A2(\sresult[19][6] ),
  .ZN(_02025_)
);

NAND2_X1 _07175_ (
  .A1(_02024_),
  .A2(_02025_),
  .ZN(_00234_)
);

NAND2_X1 _07176_ (
  .A1(_02009_),
  .A2(\sresult[18][7] ),
  .ZN(_02026_)
);

NAND2_X1 _07177_ (
  .A1(_01997_),
  .A2(din_36[7]),
  .ZN(_02027_)
);

NAND2_X1 _07178_ (
  .A1(_02026_),
  .A2(_02027_),
  .ZN(_02028_)
);

NAND2_X1 _07179_ (
  .A1(_02028_),
  .A2(_02001_),
  .ZN(_02029_)
);

NAND2_X1 _07180_ (
  .A1(_02014_),
  .A2(\sresult[19][7] ),
  .ZN(_02030_)
);

NAND2_X1 _07181_ (
  .A1(_02029_),
  .A2(_02030_),
  .ZN(_00235_)
);

NAND2_X1 _07182_ (
  .A1(_02009_),
  .A2(\sresult[18][8] ),
  .ZN(_02031_)
);

NAND2_X1 _07183_ (
  .A1(_01997_),
  .A2(din_36[8]),
  .ZN(_02032_)
);

NAND2_X1 _07184_ (
  .A1(_02031_),
  .A2(_02032_),
  .ZN(_02033_)
);

NAND2_X1 _07185_ (
  .A1(_02033_),
  .A2(_02001_),
  .ZN(_02034_)
);

NAND2_X1 _07186_ (
  .A1(_02014_),
  .A2(\sresult[19][8] ),
  .ZN(_02035_)
);

NAND2_X1 _07187_ (
  .A1(_02034_),
  .A2(_02035_),
  .ZN(_00236_)
);

NAND2_X1 _07188_ (
  .A1(_02009_),
  .A2(\sresult[18][9] ),
  .ZN(_02036_)
);

NAND2_X1 _07189_ (
  .A1(_01997_),
  .A2(din_36[9]),
  .ZN(_02037_)
);

NAND2_X1 _07190_ (
  .A1(_02036_),
  .A2(_02037_),
  .ZN(_02038_)
);

NAND2_X1 _07191_ (
  .A1(_02038_),
  .A2(_02001_),
  .ZN(_02039_)
);

NAND2_X1 _07192_ (
  .A1(_02014_),
  .A2(\sresult[19][9] ),
  .ZN(_02040_)
);

NAND2_X1 _07193_ (
  .A1(_02039_),
  .A2(_02040_),
  .ZN(_00237_)
);

NAND2_X1 _07194_ (
  .A1(_02009_),
  .A2(\sresult[18][10] ),
  .ZN(_02041_)
);

NAND2_X1 _07195_ (
  .A1(_01997_),
  .A2(din_36[10]),
  .ZN(_02042_)
);

NAND2_X1 _07196_ (
  .A1(_02041_),
  .A2(_02042_),
  .ZN(_02043_)
);

NAND2_X1 _07197_ (
  .A1(_02043_),
  .A2(_02001_),
  .ZN(_02044_)
);

NAND2_X1 _07198_ (
  .A1(_02014_),
  .A2(\sresult[19][10] ),
  .ZN(_02045_)
);

NAND2_X1 _07199_ (
  .A1(_02044_),
  .A2(_02045_),
  .ZN(_00238_)
);

NAND2_X1 _07200_ (
  .A1(_02009_),
  .A2(\sresult[18][11] ),
  .ZN(_02046_)
);

NAND2_X1 _07201_ (
  .A1(_01997_),
  .A2(din_36[11]),
  .ZN(_02047_)
);

NAND2_X1 _07202_ (
  .A1(_02046_),
  .A2(_02047_),
  .ZN(_02048_)
);

NAND2_X1 _07203_ (
  .A1(_02048_),
  .A2(_02001_),
  .ZN(_02049_)
);

NAND2_X1 _07204_ (
  .A1(_02014_),
  .A2(\sresult[19][11] ),
  .ZN(_02050_)
);

NAND2_X1 _07205_ (
  .A1(_02049_),
  .A2(_02050_),
  .ZN(_00239_)
);

NAND2_X1 _07206_ (
  .A1(_02009_),
  .A2(\sresult[19][0] ),
  .ZN(_02051_)
);

BUF_X4 _07207_ (
  .A(_01563_),
  .Z(_02052_)
);

NAND2_X1 _07208_ (
  .A1(_02052_),
  .A2(din_27[0]),
  .ZN(_02053_)
);

NAND2_X1 _07209_ (
  .A1(_02051_),
  .A2(_02053_),
  .ZN(_02054_)
);

BUF_X2 _07210_ (
  .A(_02000_),
  .Z(_02055_)
);

NAND2_X1 _07211_ (
  .A1(_02054_),
  .A2(_02055_),
  .ZN(_02056_)
);

NAND2_X1 _07212_ (
  .A1(_02014_),
  .A2(\sresult[20][0] ),
  .ZN(_02057_)
);

NAND2_X1 _07213_ (
  .A1(_02056_),
  .A2(_02057_),
  .ZN(_00240_)
);

NAND2_X1 _07214_ (
  .A1(_02009_),
  .A2(\sresult[19][1] ),
  .ZN(_02058_)
);

NAND2_X1 _07215_ (
  .A1(_02052_),
  .A2(din_27[1]),
  .ZN(_02059_)
);

NAND2_X1 _07216_ (
  .A1(_02058_),
  .A2(_02059_),
  .ZN(_02060_)
);

NAND2_X1 _07217_ (
  .A1(_02060_),
  .A2(_02055_),
  .ZN(_02061_)
);

NAND2_X1 _07218_ (
  .A1(_02014_),
  .A2(\sresult[20][1] ),
  .ZN(_02062_)
);

NAND2_X1 _07219_ (
  .A1(_02061_),
  .A2(_02062_),
  .ZN(_00241_)
);

BUF_X8 _07220_ (
  .A(_00799_),
  .Z(_02063_)
);

BUF_X4 _07221_ (
  .A(_02063_),
  .Z(_02064_)
);

NAND2_X1 _07222_ (
  .A1(_02064_),
  .A2(\sresult[19][2] ),
  .ZN(_02065_)
);

NAND2_X1 _07223_ (
  .A1(_02052_),
  .A2(din_27[2]),
  .ZN(_02066_)
);

NAND2_X1 _07224_ (
  .A1(_02065_),
  .A2(_02066_),
  .ZN(_02067_)
);

NAND2_X1 _07225_ (
  .A1(_02067_),
  .A2(_02055_),
  .ZN(_02068_)
);

BUF_X1 _07226_ (
  .A(_01580_),
  .Z(_02069_)
);

NAND2_X1 _07227_ (
  .A1(_02069_),
  .A2(\sresult[20][2] ),
  .ZN(_02070_)
);

NAND2_X1 _07228_ (
  .A1(_02068_),
  .A2(_02070_),
  .ZN(_00242_)
);

NAND2_X1 _07229_ (
  .A1(_02064_),
  .A2(\sresult[19][3] ),
  .ZN(_02071_)
);

NAND2_X1 _07230_ (
  .A1(_02052_),
  .A2(din_27[3]),
  .ZN(_02072_)
);

NAND2_X1 _07231_ (
  .A1(_02071_),
  .A2(_02072_),
  .ZN(_02073_)
);

NAND2_X1 _07232_ (
  .A1(_02073_),
  .A2(_02055_),
  .ZN(_02074_)
);

NAND2_X1 _07233_ (
  .A1(_02069_),
  .A2(\sresult[20][3] ),
  .ZN(_02075_)
);

NAND2_X1 _07234_ (
  .A1(_02074_),
  .A2(_02075_),
  .ZN(_00243_)
);

NAND2_X1 _07235_ (
  .A1(_02064_),
  .A2(\sresult[19][4] ),
  .ZN(_02076_)
);

NAND2_X1 _07236_ (
  .A1(_02052_),
  .A2(din_27[4]),
  .ZN(_02077_)
);

NAND2_X1 _07237_ (
  .A1(_02076_),
  .A2(_02077_),
  .ZN(_02078_)
);

NAND2_X1 _07238_ (
  .A1(_02078_),
  .A2(_02055_),
  .ZN(_02079_)
);

NAND2_X1 _07239_ (
  .A1(_02069_),
  .A2(\sresult[20][4] ),
  .ZN(_02080_)
);

NAND2_X1 _07240_ (
  .A1(_02079_),
  .A2(_02080_),
  .ZN(_00244_)
);

NAND2_X1 _07241_ (
  .A1(_02064_),
  .A2(\sresult[19][5] ),
  .ZN(_02081_)
);

NAND2_X1 _07242_ (
  .A1(_02052_),
  .A2(din_27[5]),
  .ZN(_02082_)
);

NAND2_X1 _07243_ (
  .A1(_02081_),
  .A2(_02082_),
  .ZN(_02083_)
);

NAND2_X1 _07244_ (
  .A1(_02083_),
  .A2(_02055_),
  .ZN(_02084_)
);

NAND2_X1 _07245_ (
  .A1(_02069_),
  .A2(\sresult[20][5] ),
  .ZN(_02085_)
);

NAND2_X1 _07246_ (
  .A1(_02084_),
  .A2(_02085_),
  .ZN(_00245_)
);

NAND2_X1 _07247_ (
  .A1(_02064_),
  .A2(\sresult[19][6] ),
  .ZN(_02086_)
);

NAND2_X1 _07248_ (
  .A1(_02052_),
  .A2(din_27[6]),
  .ZN(_02087_)
);

NAND2_X1 _07249_ (
  .A1(_02086_),
  .A2(_02087_),
  .ZN(_02088_)
);

NAND2_X1 _07250_ (
  .A1(_02088_),
  .A2(_02055_),
  .ZN(_02089_)
);

NAND2_X1 _07251_ (
  .A1(_02069_),
  .A2(\sresult[20][6] ),
  .ZN(_02090_)
);

NAND2_X1 _07252_ (
  .A1(_02089_),
  .A2(_02090_),
  .ZN(_00246_)
);

NAND2_X1 _07253_ (
  .A1(_02064_),
  .A2(\sresult[19][7] ),
  .ZN(_02091_)
);

NAND2_X1 _07254_ (
  .A1(_02052_),
  .A2(din_27[7]),
  .ZN(_02092_)
);

NAND2_X1 _07255_ (
  .A1(_02091_),
  .A2(_02092_),
  .ZN(_02093_)
);

NAND2_X1 _07256_ (
  .A1(_02093_),
  .A2(_02055_),
  .ZN(_02094_)
);

NAND2_X1 _07257_ (
  .A1(_02069_),
  .A2(\sresult[20][7] ),
  .ZN(_02095_)
);

NAND2_X1 _07258_ (
  .A1(_02094_),
  .A2(_02095_),
  .ZN(_00247_)
);

NAND2_X1 _07259_ (
  .A1(_02064_),
  .A2(\sresult[19][8] ),
  .ZN(_02096_)
);

NAND2_X1 _07260_ (
  .A1(_02052_),
  .A2(din_27[8]),
  .ZN(_02097_)
);

NAND2_X1 _07261_ (
  .A1(_02096_),
  .A2(_02097_),
  .ZN(_02098_)
);

NAND2_X1 _07262_ (
  .A1(_02098_),
  .A2(_02055_),
  .ZN(_02099_)
);

NAND2_X1 _07263_ (
  .A1(_02069_),
  .A2(\sresult[20][8] ),
  .ZN(_02100_)
);

NAND2_X1 _07264_ (
  .A1(_02099_),
  .A2(_02100_),
  .ZN(_00248_)
);

NAND2_X1 _07265_ (
  .A1(_02064_),
  .A2(\sresult[19][9] ),
  .ZN(_02101_)
);

NAND2_X1 _07266_ (
  .A1(_02052_),
  .A2(din_27[9]),
  .ZN(_02102_)
);

NAND2_X1 _07267_ (
  .A1(_02101_),
  .A2(_02102_),
  .ZN(_02103_)
);

NAND2_X1 _07268_ (
  .A1(_02103_),
  .A2(_02055_),
  .ZN(_02104_)
);

NAND2_X1 _07269_ (
  .A1(_02069_),
  .A2(\sresult[20][9] ),
  .ZN(_02105_)
);

NAND2_X1 _07270_ (
  .A1(_02104_),
  .A2(_02105_),
  .ZN(_00249_)
);

NAND2_X1 _07271_ (
  .A1(_02064_),
  .A2(\sresult[19][10] ),
  .ZN(_02106_)
);

BUF_X8 _07272_ (
  .A(_00770_),
  .Z(_02107_)
);

BUF_X4 _07273_ (
  .A(_02107_),
  .Z(_02108_)
);

NAND2_X1 _07274_ (
  .A1(_02108_),
  .A2(din_27[10]),
  .ZN(_02109_)
);

NAND2_X1 _07275_ (
  .A1(_02106_),
  .A2(_02109_),
  .ZN(_02110_)
);

BUF_X2 _07276_ (
  .A(_02000_),
  .Z(_02111_)
);

NAND2_X1 _07277_ (
  .A1(_02110_),
  .A2(_02111_),
  .ZN(_02112_)
);

NAND2_X1 _07278_ (
  .A1(_02069_),
  .A2(\sresult[20][10] ),
  .ZN(_02113_)
);

NAND2_X1 _07279_ (
  .A1(_02112_),
  .A2(_02113_),
  .ZN(_00250_)
);

NAND2_X1 _07280_ (
  .A1(_02064_),
  .A2(\sresult[19][11] ),
  .ZN(_02114_)
);

NAND2_X1 _07281_ (
  .A1(_02108_),
  .A2(din_27[11]),
  .ZN(_02115_)
);

NAND2_X1 _07282_ (
  .A1(_02114_),
  .A2(_02115_),
  .ZN(_02116_)
);

NAND2_X1 _07283_ (
  .A1(_02116_),
  .A2(_02111_),
  .ZN(_02117_)
);

NAND2_X1 _07284_ (
  .A1(_02069_),
  .A2(\sresult[20][11] ),
  .ZN(_02118_)
);

NAND2_X1 _07285_ (
  .A1(_02117_),
  .A2(_02118_),
  .ZN(_00251_)
);

BUF_X4 _07286_ (
  .A(_02063_),
  .Z(_02119_)
);

NAND2_X1 _07287_ (
  .A1(_02119_),
  .A2(\sresult[20][0] ),
  .ZN(_02120_)
);

NAND2_X1 _07288_ (
  .A1(_02108_),
  .A2(din_17[0]),
  .ZN(_02121_)
);

NAND2_X1 _07289_ (
  .A1(_02120_),
  .A2(_02121_),
  .ZN(_02122_)
);

NAND2_X1 _07290_ (
  .A1(_02122_),
  .A2(_02111_),
  .ZN(_02123_)
);

BUF_X8 _07291_ (
  .A(_00810_),
  .Z(_02124_)
);

BUF_X1 _07292_ (
  .A(_02124_),
  .Z(_02125_)
);

NAND2_X1 _07293_ (
  .A1(_02125_),
  .A2(\sresult[21][0] ),
  .ZN(_02126_)
);

NAND2_X1 _07294_ (
  .A1(_02123_),
  .A2(_02126_),
  .ZN(_00252_)
);

NAND2_X1 _07295_ (
  .A1(_02119_),
  .A2(\sresult[20][1] ),
  .ZN(_02127_)
);

NAND2_X1 _07296_ (
  .A1(_02108_),
  .A2(din_17[1]),
  .ZN(_02128_)
);

NAND2_X1 _07297_ (
  .A1(_02127_),
  .A2(_02128_),
  .ZN(_02129_)
);

NAND2_X1 _07298_ (
  .A1(_02129_),
  .A2(_02111_),
  .ZN(_02130_)
);

NAND2_X1 _07299_ (
  .A1(_02125_),
  .A2(\sresult[21][1] ),
  .ZN(_02131_)
);

NAND2_X1 _07300_ (
  .A1(_02130_),
  .A2(_02131_),
  .ZN(_00253_)
);

NAND2_X1 _07301_ (
  .A1(_02119_),
  .A2(\sresult[20][2] ),
  .ZN(_02132_)
);

NAND2_X1 _07302_ (
  .A1(_02108_),
  .A2(din_17[2]),
  .ZN(_02133_)
);

NAND2_X1 _07303_ (
  .A1(_02132_),
  .A2(_02133_),
  .ZN(_02134_)
);

NAND2_X1 _07304_ (
  .A1(_02134_),
  .A2(_02111_),
  .ZN(_02135_)
);

NAND2_X1 _07305_ (
  .A1(_02125_),
  .A2(\sresult[21][2] ),
  .ZN(_02136_)
);

NAND2_X1 _07306_ (
  .A1(_02135_),
  .A2(_02136_),
  .ZN(_00254_)
);

NAND2_X1 _07307_ (
  .A1(_02119_),
  .A2(\sresult[20][3] ),
  .ZN(_02137_)
);

NAND2_X1 _07308_ (
  .A1(_02108_),
  .A2(din_17[3]),
  .ZN(_02138_)
);

NAND2_X1 _07309_ (
  .A1(_02137_),
  .A2(_02138_),
  .ZN(_02139_)
);

NAND2_X1 _07310_ (
  .A1(_02139_),
  .A2(_02111_),
  .ZN(_02140_)
);

NAND2_X1 _07311_ (
  .A1(_02125_),
  .A2(\sresult[21][3] ),
  .ZN(_02141_)
);

NAND2_X1 _07312_ (
  .A1(_02140_),
  .A2(_02141_),
  .ZN(_00255_)
);

NAND2_X1 _07313_ (
  .A1(_02119_),
  .A2(\sresult[20][4] ),
  .ZN(_02142_)
);

NAND2_X1 _07314_ (
  .A1(_02108_),
  .A2(din_17[4]),
  .ZN(_02143_)
);

NAND2_X1 _07315_ (
  .A1(_02142_),
  .A2(_02143_),
  .ZN(_02144_)
);

NAND2_X1 _07316_ (
  .A1(_02144_),
  .A2(_02111_),
  .ZN(_02145_)
);

NAND2_X1 _07317_ (
  .A1(_02125_),
  .A2(\sresult[21][4] ),
  .ZN(_02146_)
);

NAND2_X1 _07318_ (
  .A1(_02145_),
  .A2(_02146_),
  .ZN(_00256_)
);

NAND2_X1 _07319_ (
  .A1(_02119_),
  .A2(\sresult[20][5] ),
  .ZN(_02147_)
);

NAND2_X1 _07320_ (
  .A1(_02108_),
  .A2(din_17[5]),
  .ZN(_02148_)
);

NAND2_X1 _07321_ (
  .A1(_02147_),
  .A2(_02148_),
  .ZN(_02149_)
);

NAND2_X1 _07322_ (
  .A1(_02149_),
  .A2(_02111_),
  .ZN(_02150_)
);

NAND2_X1 _07323_ (
  .A1(_02125_),
  .A2(\sresult[21][5] ),
  .ZN(_02151_)
);

NAND2_X1 _07324_ (
  .A1(_02150_),
  .A2(_02151_),
  .ZN(_00257_)
);

NAND2_X1 _07325_ (
  .A1(_02119_),
  .A2(\sresult[20][6] ),
  .ZN(_02152_)
);

NAND2_X1 _07326_ (
  .A1(_02108_),
  .A2(din_17[6]),
  .ZN(_02153_)
);

NAND2_X1 _07327_ (
  .A1(_02152_),
  .A2(_02153_),
  .ZN(_02154_)
);

NAND2_X1 _07328_ (
  .A1(_02154_),
  .A2(_02111_),
  .ZN(_02155_)
);

NAND2_X1 _07329_ (
  .A1(_02125_),
  .A2(\sresult[21][6] ),
  .ZN(_02156_)
);

NAND2_X1 _07330_ (
  .A1(_02155_),
  .A2(_02156_),
  .ZN(_00258_)
);

NAND2_X1 _07331_ (
  .A1(_02119_),
  .A2(\sresult[20][7] ),
  .ZN(_02157_)
);

NAND2_X1 _07332_ (
  .A1(_02108_),
  .A2(din_17[7]),
  .ZN(_02158_)
);

NAND2_X1 _07333_ (
  .A1(_02157_),
  .A2(_02158_),
  .ZN(_02159_)
);

NAND2_X1 _07334_ (
  .A1(_02159_),
  .A2(_02111_),
  .ZN(_02160_)
);

NAND2_X1 _07335_ (
  .A1(_02125_),
  .A2(\sresult[21][7] ),
  .ZN(_02161_)
);

NAND2_X1 _07336_ (
  .A1(_02160_),
  .A2(_02161_),
  .ZN(_00259_)
);

NAND2_X1 _07337_ (
  .A1(_02119_),
  .A2(\sresult[20][8] ),
  .ZN(_02162_)
);

BUF_X4 _07338_ (
  .A(_02107_),
  .Z(_02163_)
);

NAND2_X1 _07339_ (
  .A1(_02163_),
  .A2(din_17[8]),
  .ZN(_02164_)
);

NAND2_X1 _07340_ (
  .A1(_02162_),
  .A2(_02164_),
  .ZN(_02165_)
);

BUF_X2 _07341_ (
  .A(_02000_),
  .Z(_02166_)
);

NAND2_X1 _07342_ (
  .A1(_02165_),
  .A2(_02166_),
  .ZN(_02167_)
);

NAND2_X1 _07343_ (
  .A1(_02125_),
  .A2(\sresult[21][8] ),
  .ZN(_02168_)
);

NAND2_X1 _07344_ (
  .A1(_02167_),
  .A2(_02168_),
  .ZN(_00260_)
);

NAND2_X1 _07345_ (
  .A1(_02119_),
  .A2(\sresult[20][9] ),
  .ZN(_02169_)
);

NAND2_X1 _07346_ (
  .A1(_02163_),
  .A2(din_17[9]),
  .ZN(_02170_)
);

NAND2_X1 _07347_ (
  .A1(_02169_),
  .A2(_02170_),
  .ZN(_02171_)
);

NAND2_X1 _07348_ (
  .A1(_02171_),
  .A2(_02166_),
  .ZN(_02172_)
);

NAND2_X1 _07349_ (
  .A1(_02125_),
  .A2(\sresult[21][9] ),
  .ZN(_02173_)
);

NAND2_X1 _07350_ (
  .A1(_02172_),
  .A2(_02173_),
  .ZN(_00261_)
);

BUF_X4 _07351_ (
  .A(_02063_),
  .Z(_02174_)
);

NAND2_X1 _07352_ (
  .A1(_02174_),
  .A2(\sresult[20][10] ),
  .ZN(_02175_)
);

NAND2_X1 _07353_ (
  .A1(_02163_),
  .A2(din_17[10]),
  .ZN(_02176_)
);

NAND2_X1 _07354_ (
  .A1(_02175_),
  .A2(_02176_),
  .ZN(_02177_)
);

NAND2_X1 _07355_ (
  .A1(_02177_),
  .A2(_02166_),
  .ZN(_02178_)
);

BUF_X1 _07356_ (
  .A(_02124_),
  .Z(_02179_)
);

NAND2_X1 _07357_ (
  .A1(_02179_),
  .A2(\sresult[21][10] ),
  .ZN(_02180_)
);

NAND2_X1 _07358_ (
  .A1(_02178_),
  .A2(_02180_),
  .ZN(_00262_)
);

NAND2_X1 _07359_ (
  .A1(_02174_),
  .A2(\sresult[20][11] ),
  .ZN(_02181_)
);

NAND2_X1 _07360_ (
  .A1(_02163_),
  .A2(din_17[11]),
  .ZN(_02182_)
);

NAND2_X1 _07361_ (
  .A1(_02181_),
  .A2(_02182_),
  .ZN(_02183_)
);

NAND2_X1 _07362_ (
  .A1(_02183_),
  .A2(_02166_),
  .ZN(_02184_)
);

NAND2_X1 _07363_ (
  .A1(_02179_),
  .A2(\sresult[21][11] ),
  .ZN(_02185_)
);

NAND2_X1 _07364_ (
  .A1(_02184_),
  .A2(_02185_),
  .ZN(_00263_)
);

NAND2_X1 _07365_ (
  .A1(_02174_),
  .A2(\sresult[21][0] ),
  .ZN(_02186_)
);

NAND2_X1 _07366_ (
  .A1(_02163_),
  .A2(din_26[0]),
  .ZN(_02187_)
);

NAND2_X1 _07367_ (
  .A1(_02186_),
  .A2(_02187_),
  .ZN(_02188_)
);

NAND2_X1 _07368_ (
  .A1(_02188_),
  .A2(_02166_),
  .ZN(_02189_)
);

NAND2_X1 _07369_ (
  .A1(_02179_),
  .A2(\sresult[22][0] ),
  .ZN(_02190_)
);

NAND2_X1 _07370_ (
  .A1(_02189_),
  .A2(_02190_),
  .ZN(_00264_)
);

NAND2_X1 _07371_ (
  .A1(_02174_),
  .A2(\sresult[21][1] ),
  .ZN(_02191_)
);

NAND2_X1 _07372_ (
  .A1(_02163_),
  .A2(din_26[1]),
  .ZN(_02192_)
);

NAND2_X1 _07373_ (
  .A1(_02191_),
  .A2(_02192_),
  .ZN(_02193_)
);

NAND2_X1 _07374_ (
  .A1(_02193_),
  .A2(_02166_),
  .ZN(_02194_)
);

NAND2_X1 _07375_ (
  .A1(_02179_),
  .A2(\sresult[22][1] ),
  .ZN(_02195_)
);

NAND2_X1 _07376_ (
  .A1(_02194_),
  .A2(_02195_),
  .ZN(_00265_)
);

NAND2_X1 _07377_ (
  .A1(_02174_),
  .A2(\sresult[21][2] ),
  .ZN(_02196_)
);

NAND2_X1 _07378_ (
  .A1(_02163_),
  .A2(din_26[2]),
  .ZN(_02197_)
);

NAND2_X1 _07379_ (
  .A1(_02196_),
  .A2(_02197_),
  .ZN(_02198_)
);

NAND2_X1 _07380_ (
  .A1(_02198_),
  .A2(_02166_),
  .ZN(_02199_)
);

NAND2_X1 _07381_ (
  .A1(_02179_),
  .A2(\sresult[22][2] ),
  .ZN(_02200_)
);

NAND2_X1 _07382_ (
  .A1(_02199_),
  .A2(_02200_),
  .ZN(_00266_)
);

NAND2_X1 _07383_ (
  .A1(_02174_),
  .A2(\sresult[21][3] ),
  .ZN(_02201_)
);

NAND2_X1 _07384_ (
  .A1(_02163_),
  .A2(din_26[3]),
  .ZN(_02202_)
);

NAND2_X1 _07385_ (
  .A1(_02201_),
  .A2(_02202_),
  .ZN(_02203_)
);

NAND2_X1 _07386_ (
  .A1(_02203_),
  .A2(_02166_),
  .ZN(_02204_)
);

NAND2_X1 _07387_ (
  .A1(_02179_),
  .A2(\sresult[22][3] ),
  .ZN(_02205_)
);

NAND2_X1 _07388_ (
  .A1(_02204_),
  .A2(_02205_),
  .ZN(_00267_)
);

NAND2_X1 _07389_ (
  .A1(_02174_),
  .A2(\sresult[21][4] ),
  .ZN(_02206_)
);

NAND2_X1 _07390_ (
  .A1(_02163_),
  .A2(din_26[4]),
  .ZN(_02207_)
);

NAND2_X1 _07391_ (
  .A1(_02206_),
  .A2(_02207_),
  .ZN(_02208_)
);

NAND2_X1 _07392_ (
  .A1(_02208_),
  .A2(_02166_),
  .ZN(_02209_)
);

NAND2_X1 _07393_ (
  .A1(_02179_),
  .A2(\sresult[22][4] ),
  .ZN(_02210_)
);

NAND2_X1 _07394_ (
  .A1(_02209_),
  .A2(_02210_),
  .ZN(_00268_)
);

NAND2_X1 _07395_ (
  .A1(_02174_),
  .A2(\sresult[21][5] ),
  .ZN(_02211_)
);

NAND2_X1 _07396_ (
  .A1(_02163_),
  .A2(din_26[5]),
  .ZN(_02212_)
);

NAND2_X1 _07397_ (
  .A1(_02211_),
  .A2(_02212_),
  .ZN(_02213_)
);

NAND2_X1 _07398_ (
  .A1(_02213_),
  .A2(_02166_),
  .ZN(_02214_)
);

NAND2_X1 _07399_ (
  .A1(_02179_),
  .A2(\sresult[22][5] ),
  .ZN(_02215_)
);

NAND2_X1 _07400_ (
  .A1(_02214_),
  .A2(_02215_),
  .ZN(_00269_)
);

NAND2_X1 _07401_ (
  .A1(_02174_),
  .A2(\sresult[21][6] ),
  .ZN(_02216_)
);

BUF_X4 _07402_ (
  .A(_02107_),
  .Z(_02217_)
);

NAND2_X1 _07403_ (
  .A1(_02217_),
  .A2(din_26[6]),
  .ZN(_02218_)
);

NAND2_X1 _07404_ (
  .A1(_02216_),
  .A2(_02218_),
  .ZN(_02219_)
);

BUF_X2 _07405_ (
  .A(_02000_),
  .Z(_02220_)
);

NAND2_X1 _07406_ (
  .A1(_02219_),
  .A2(_02220_),
  .ZN(_02221_)
);

NAND2_X1 _07407_ (
  .A1(_02179_),
  .A2(\sresult[22][6] ),
  .ZN(_02222_)
);

NAND2_X1 _07408_ (
  .A1(_02221_),
  .A2(_02222_),
  .ZN(_00270_)
);

NAND2_X1 _07409_ (
  .A1(_02174_),
  .A2(\sresult[21][7] ),
  .ZN(_02223_)
);

NAND2_X1 _07410_ (
  .A1(_02217_),
  .A2(din_26[7]),
  .ZN(_02224_)
);

NAND2_X1 _07411_ (
  .A1(_02223_),
  .A2(_02224_),
  .ZN(_02225_)
);

NAND2_X1 _07412_ (
  .A1(_02225_),
  .A2(_02220_),
  .ZN(_02226_)
);

NAND2_X1 _07413_ (
  .A1(_02179_),
  .A2(\sresult[22][7] ),
  .ZN(_02227_)
);

NAND2_X1 _07414_ (
  .A1(_02226_),
  .A2(_02227_),
  .ZN(_00271_)
);

BUF_X4 _07415_ (
  .A(_02063_),
  .Z(_02228_)
);

NAND2_X1 _07416_ (
  .A1(_02228_),
  .A2(\sresult[21][8] ),
  .ZN(_02229_)
);

NAND2_X1 _07417_ (
  .A1(_02217_),
  .A2(din_26[8]),
  .ZN(_02230_)
);

NAND2_X1 _07418_ (
  .A1(_02229_),
  .A2(_02230_),
  .ZN(_02231_)
);

NAND2_X1 _07419_ (
  .A1(_02231_),
  .A2(_02220_),
  .ZN(_02232_)
);

BUF_X1 _07420_ (
  .A(_02124_),
  .Z(_02233_)
);

NAND2_X1 _07421_ (
  .A1(_02233_),
  .A2(\sresult[22][8] ),
  .ZN(_02234_)
);

NAND2_X1 _07422_ (
  .A1(_02232_),
  .A2(_02234_),
  .ZN(_00272_)
);

NAND2_X1 _07423_ (
  .A1(_02228_),
  .A2(\sresult[21][9] ),
  .ZN(_02235_)
);

NAND2_X1 _07424_ (
  .A1(_02217_),
  .A2(din_26[9]),
  .ZN(_02236_)
);

NAND2_X1 _07425_ (
  .A1(_02235_),
  .A2(_02236_),
  .ZN(_02237_)
);

NAND2_X1 _07426_ (
  .A1(_02237_),
  .A2(_02220_),
  .ZN(_02238_)
);

NAND2_X1 _07427_ (
  .A1(_02233_),
  .A2(\sresult[22][9] ),
  .ZN(_02239_)
);

NAND2_X1 _07428_ (
  .A1(_02238_),
  .A2(_02239_),
  .ZN(_00273_)
);

NAND2_X1 _07429_ (
  .A1(_02228_),
  .A2(\sresult[21][10] ),
  .ZN(_02240_)
);

NAND2_X1 _07430_ (
  .A1(_02217_),
  .A2(din_26[10]),
  .ZN(_02241_)
);

NAND2_X1 _07431_ (
  .A1(_02240_),
  .A2(_02241_),
  .ZN(_02242_)
);

NAND2_X1 _07432_ (
  .A1(_02242_),
  .A2(_02220_),
  .ZN(_02243_)
);

NAND2_X1 _07433_ (
  .A1(_02233_),
  .A2(\sresult[22][10] ),
  .ZN(_02244_)
);

NAND2_X1 _07434_ (
  .A1(_02243_),
  .A2(_02244_),
  .ZN(_00274_)
);

NAND2_X1 _07435_ (
  .A1(_02228_),
  .A2(\sresult[21][11] ),
  .ZN(_02245_)
);

NAND2_X1 _07436_ (
  .A1(_02217_),
  .A2(din_26[11]),
  .ZN(_02246_)
);

NAND2_X1 _07437_ (
  .A1(_02245_),
  .A2(_02246_),
  .ZN(_02247_)
);

NAND2_X1 _07438_ (
  .A1(_02247_),
  .A2(_02220_),
  .ZN(_02248_)
);

NAND2_X1 _07439_ (
  .A1(_02233_),
  .A2(\sresult[22][11] ),
  .ZN(_02249_)
);

NAND2_X1 _07440_ (
  .A1(_02248_),
  .A2(_02249_),
  .ZN(_00275_)
);

NAND2_X1 _07441_ (
  .A1(_02228_),
  .A2(\sresult[22][0] ),
  .ZN(_02250_)
);

NAND2_X1 _07442_ (
  .A1(_02217_),
  .A2(din_35[0]),
  .ZN(_02251_)
);

NAND2_X1 _07443_ (
  .A1(_02250_),
  .A2(_02251_),
  .ZN(_02252_)
);

NAND2_X1 _07444_ (
  .A1(_02252_),
  .A2(_02220_),
  .ZN(_02253_)
);

NAND2_X1 _07445_ (
  .A1(_02233_),
  .A2(\sresult[23][0] ),
  .ZN(_02254_)
);

NAND2_X1 _07446_ (
  .A1(_02253_),
  .A2(_02254_),
  .ZN(_00276_)
);

NAND2_X1 _07447_ (
  .A1(_02228_),
  .A2(\sresult[22][1] ),
  .ZN(_02255_)
);

NAND2_X1 _07448_ (
  .A1(_02217_),
  .A2(din_35[1]),
  .ZN(_02256_)
);

NAND2_X1 _07449_ (
  .A1(_02255_),
  .A2(_02256_),
  .ZN(_02257_)
);

NAND2_X1 _07450_ (
  .A1(_02257_),
  .A2(_02220_),
  .ZN(_02258_)
);

NAND2_X1 _07451_ (
  .A1(_02233_),
  .A2(\sresult[23][1] ),
  .ZN(_02259_)
);

NAND2_X1 _07452_ (
  .A1(_02258_),
  .A2(_02259_),
  .ZN(_00277_)
);

NAND2_X1 _07453_ (
  .A1(_02228_),
  .A2(\sresult[22][2] ),
  .ZN(_02260_)
);

NAND2_X1 _07454_ (
  .A1(_02217_),
  .A2(din_35[2]),
  .ZN(_02261_)
);

NAND2_X1 _07455_ (
  .A1(_02260_),
  .A2(_02261_),
  .ZN(_02262_)
);

NAND2_X1 _07456_ (
  .A1(_02262_),
  .A2(_02220_),
  .ZN(_02263_)
);

NAND2_X1 _07457_ (
  .A1(_02233_),
  .A2(\sresult[23][2] ),
  .ZN(_02264_)
);

NAND2_X1 _07458_ (
  .A1(_02263_),
  .A2(_02264_),
  .ZN(_00278_)
);

NAND2_X1 _07459_ (
  .A1(_02228_),
  .A2(\sresult[22][3] ),
  .ZN(_02265_)
);

NAND2_X1 _07460_ (
  .A1(_02217_),
  .A2(din_35[3]),
  .ZN(_02266_)
);

NAND2_X1 _07461_ (
  .A1(_02265_),
  .A2(_02266_),
  .ZN(_02267_)
);

NAND2_X1 _07462_ (
  .A1(_02267_),
  .A2(_02220_),
  .ZN(_02268_)
);

NAND2_X1 _07463_ (
  .A1(_02233_),
  .A2(\sresult[23][3] ),
  .ZN(_02269_)
);

NAND2_X1 _07464_ (
  .A1(_02268_),
  .A2(_02269_),
  .ZN(_00279_)
);

NAND2_X1 _07465_ (
  .A1(_02228_),
  .A2(\sresult[22][4] ),
  .ZN(_02270_)
);

BUF_X4 _07466_ (
  .A(_02107_),
  .Z(_02271_)
);

NAND2_X1 _07467_ (
  .A1(_02271_),
  .A2(din_35[4]),
  .ZN(_02272_)
);

NAND2_X1 _07468_ (
  .A1(_02270_),
  .A2(_02272_),
  .ZN(_02273_)
);

BUF_X2 _07469_ (
  .A(_02000_),
  .Z(_02274_)
);

NAND2_X1 _07470_ (
  .A1(_02273_),
  .A2(_02274_),
  .ZN(_02275_)
);

NAND2_X1 _07471_ (
  .A1(_02233_),
  .A2(\sresult[23][4] ),
  .ZN(_02276_)
);

NAND2_X1 _07472_ (
  .A1(_02275_),
  .A2(_02276_),
  .ZN(_00280_)
);

NAND2_X1 _07473_ (
  .A1(_02228_),
  .A2(\sresult[22][5] ),
  .ZN(_02277_)
);

NAND2_X1 _07474_ (
  .A1(_02271_),
  .A2(din_35[5]),
  .ZN(_02278_)
);

NAND2_X1 _07475_ (
  .A1(_02277_),
  .A2(_02278_),
  .ZN(_02279_)
);

NAND2_X1 _07476_ (
  .A1(_02279_),
  .A2(_02274_),
  .ZN(_02280_)
);

NAND2_X1 _07477_ (
  .A1(_02233_),
  .A2(\sresult[23][5] ),
  .ZN(_02281_)
);

NAND2_X1 _07478_ (
  .A1(_02280_),
  .A2(_02281_),
  .ZN(_00281_)
);

BUF_X4 _07479_ (
  .A(_02063_),
  .Z(_02282_)
);

NAND2_X1 _07480_ (
  .A1(_02282_),
  .A2(\sresult[22][6] ),
  .ZN(_02283_)
);

NAND2_X1 _07481_ (
  .A1(_02271_),
  .A2(din_35[6]),
  .ZN(_02284_)
);

NAND2_X1 _07482_ (
  .A1(_02283_),
  .A2(_02284_),
  .ZN(_02285_)
);

NAND2_X1 _07483_ (
  .A1(_02285_),
  .A2(_02274_),
  .ZN(_02286_)
);

BUF_X1 _07484_ (
  .A(_02124_),
  .Z(_02287_)
);

NAND2_X1 _07485_ (
  .A1(_02287_),
  .A2(\sresult[23][6] ),
  .ZN(_02288_)
);

NAND2_X1 _07486_ (
  .A1(_02286_),
  .A2(_02288_),
  .ZN(_00282_)
);

NAND2_X1 _07487_ (
  .A1(_02282_),
  .A2(\sresult[22][7] ),
  .ZN(_02289_)
);

NAND2_X1 _07488_ (
  .A1(_02271_),
  .A2(din_35[7]),
  .ZN(_02290_)
);

NAND2_X1 _07489_ (
  .A1(_02289_),
  .A2(_02290_),
  .ZN(_02291_)
);

NAND2_X1 _07490_ (
  .A1(_02291_),
  .A2(_02274_),
  .ZN(_02292_)
);

NAND2_X1 _07491_ (
  .A1(_02287_),
  .A2(\sresult[23][7] ),
  .ZN(_02293_)
);

NAND2_X1 _07492_ (
  .A1(_02292_),
  .A2(_02293_),
  .ZN(_00283_)
);

NAND2_X1 _07493_ (
  .A1(_02282_),
  .A2(\sresult[22][8] ),
  .ZN(_02294_)
);

NAND2_X1 _07494_ (
  .A1(_02271_),
  .A2(din_35[8]),
  .ZN(_02295_)
);

NAND2_X1 _07495_ (
  .A1(_02294_),
  .A2(_02295_),
  .ZN(_02296_)
);

NAND2_X1 _07496_ (
  .A1(_02296_),
  .A2(_02274_),
  .ZN(_02297_)
);

NAND2_X1 _07497_ (
  .A1(_02287_),
  .A2(\sresult[23][8] ),
  .ZN(_02298_)
);

NAND2_X1 _07498_ (
  .A1(_02297_),
  .A2(_02298_),
  .ZN(_00284_)
);

NAND2_X1 _07499_ (
  .A1(_02282_),
  .A2(\sresult[22][9] ),
  .ZN(_02299_)
);

NAND2_X1 _07500_ (
  .A1(_02271_),
  .A2(din_35[9]),
  .ZN(_02300_)
);

NAND2_X1 _07501_ (
  .A1(_02299_),
  .A2(_02300_),
  .ZN(_02301_)
);

NAND2_X1 _07502_ (
  .A1(_02301_),
  .A2(_02274_),
  .ZN(_02302_)
);

NAND2_X1 _07503_ (
  .A1(_02287_),
  .A2(\sresult[23][9] ),
  .ZN(_02303_)
);

NAND2_X1 _07504_ (
  .A1(_02302_),
  .A2(_02303_),
  .ZN(_00285_)
);

NAND2_X1 _07505_ (
  .A1(_02282_),
  .A2(\sresult[22][10] ),
  .ZN(_02304_)
);

NAND2_X1 _07506_ (
  .A1(_02271_),
  .A2(din_35[10]),
  .ZN(_02305_)
);

NAND2_X1 _07507_ (
  .A1(_02304_),
  .A2(_02305_),
  .ZN(_02306_)
);

NAND2_X1 _07508_ (
  .A1(_02306_),
  .A2(_02274_),
  .ZN(_02307_)
);

NAND2_X1 _07509_ (
  .A1(_02287_),
  .A2(\sresult[23][10] ),
  .ZN(_02308_)
);

NAND2_X1 _07510_ (
  .A1(_02307_),
  .A2(_02308_),
  .ZN(_00286_)
);

NAND2_X1 _07511_ (
  .A1(_02282_),
  .A2(\sresult[22][11] ),
  .ZN(_02309_)
);

NAND2_X1 _07512_ (
  .A1(_02271_),
  .A2(din_35[11]),
  .ZN(_02310_)
);

NAND2_X1 _07513_ (
  .A1(_02309_),
  .A2(_02310_),
  .ZN(_02311_)
);

NAND2_X1 _07514_ (
  .A1(_02311_),
  .A2(_02274_),
  .ZN(_02312_)
);

NAND2_X1 _07515_ (
  .A1(_02287_),
  .A2(\sresult[23][11] ),
  .ZN(_02313_)
);

NAND2_X1 _07516_ (
  .A1(_02312_),
  .A2(_02313_),
  .ZN(_00287_)
);

NAND2_X1 _07517_ (
  .A1(_02282_),
  .A2(\sresult[23][0] ),
  .ZN(_02314_)
);

NAND2_X1 _07518_ (
  .A1(_02271_),
  .A2(din_44[0]),
  .ZN(_02315_)
);

NAND2_X1 _07519_ (
  .A1(_02314_),
  .A2(_02315_),
  .ZN(_02316_)
);

NAND2_X1 _07520_ (
  .A1(_02316_),
  .A2(_02274_),
  .ZN(_02317_)
);

NAND2_X1 _07521_ (
  .A1(_02287_),
  .A2(\sresult[24][0] ),
  .ZN(_02318_)
);

NAND2_X1 _07522_ (
  .A1(_02317_),
  .A2(_02318_),
  .ZN(_00288_)
);

NAND2_X1 _07523_ (
  .A1(_02282_),
  .A2(\sresult[23][1] ),
  .ZN(_02319_)
);

NAND2_X1 _07524_ (
  .A1(_02271_),
  .A2(din_44[1]),
  .ZN(_02320_)
);

NAND2_X1 _07525_ (
  .A1(_02319_),
  .A2(_02320_),
  .ZN(_02321_)
);

NAND2_X1 _07526_ (
  .A1(_02321_),
  .A2(_02274_),
  .ZN(_02322_)
);

NAND2_X1 _07527_ (
  .A1(_02287_),
  .A2(\sresult[24][1] ),
  .ZN(_02323_)
);

NAND2_X1 _07528_ (
  .A1(_02322_),
  .A2(_02323_),
  .ZN(_00289_)
);

NAND2_X1 _07529_ (
  .A1(_02282_),
  .A2(\sresult[23][2] ),
  .ZN(_02324_)
);

BUF_X4 _07530_ (
  .A(_02107_),
  .Z(_02325_)
);

NAND2_X1 _07531_ (
  .A1(_02325_),
  .A2(din_44[2]),
  .ZN(_02326_)
);

NAND2_X1 _07532_ (
  .A1(_02324_),
  .A2(_02326_),
  .ZN(_02327_)
);

BUF_X2 _07533_ (
  .A(_02000_),
  .Z(_02328_)
);

NAND2_X1 _07534_ (
  .A1(_02327_),
  .A2(_02328_),
  .ZN(_02329_)
);

NAND2_X1 _07535_ (
  .A1(_02287_),
  .A2(\sresult[24][2] ),
  .ZN(_02330_)
);

NAND2_X1 _07536_ (
  .A1(_02329_),
  .A2(_02330_),
  .ZN(_00290_)
);

NAND2_X1 _07537_ (
  .A1(_02282_),
  .A2(\sresult[23][3] ),
  .ZN(_02331_)
);

NAND2_X1 _07538_ (
  .A1(_02325_),
  .A2(din_44[3]),
  .ZN(_02332_)
);

NAND2_X1 _07539_ (
  .A1(_02331_),
  .A2(_02332_),
  .ZN(_02333_)
);

NAND2_X1 _07540_ (
  .A1(_02333_),
  .A2(_02328_),
  .ZN(_02334_)
);

NAND2_X1 _07541_ (
  .A1(_02287_),
  .A2(\sresult[24][3] ),
  .ZN(_02335_)
);

NAND2_X1 _07542_ (
  .A1(_02334_),
  .A2(_02335_),
  .ZN(_00291_)
);

BUF_X4 _07543_ (
  .A(_02063_),
  .Z(_02336_)
);

NAND2_X1 _07544_ (
  .A1(_02336_),
  .A2(\sresult[23][4] ),
  .ZN(_02337_)
);

NAND2_X1 _07545_ (
  .A1(_02325_),
  .A2(din_44[4]),
  .ZN(_02338_)
);

NAND2_X1 _07546_ (
  .A1(_02337_),
  .A2(_02338_),
  .ZN(_02339_)
);

NAND2_X1 _07547_ (
  .A1(_02339_),
  .A2(_02328_),
  .ZN(_02340_)
);

BUF_X1 _07548_ (
  .A(_02124_),
  .Z(_02341_)
);

NAND2_X1 _07549_ (
  .A1(_02341_),
  .A2(\sresult[24][4] ),
  .ZN(_02342_)
);

NAND2_X1 _07550_ (
  .A1(_02340_),
  .A2(_02342_),
  .ZN(_00292_)
);

NAND2_X1 _07551_ (
  .A1(_02336_),
  .A2(\sresult[23][5] ),
  .ZN(_02343_)
);

NAND2_X1 _07552_ (
  .A1(_02325_),
  .A2(din_44[5]),
  .ZN(_02344_)
);

NAND2_X1 _07553_ (
  .A1(_02343_),
  .A2(_02344_),
  .ZN(_02345_)
);

NAND2_X1 _07554_ (
  .A1(_02345_),
  .A2(_02328_),
  .ZN(_02346_)
);

NAND2_X1 _07555_ (
  .A1(_02341_),
  .A2(\sresult[24][5] ),
  .ZN(_02347_)
);

NAND2_X1 _07556_ (
  .A1(_02346_),
  .A2(_02347_),
  .ZN(_00293_)
);

NAND2_X1 _07557_ (
  .A1(_02336_),
  .A2(\sresult[23][6] ),
  .ZN(_02348_)
);

NAND2_X1 _07558_ (
  .A1(_02325_),
  .A2(din_44[6]),
  .ZN(_02349_)
);

NAND2_X1 _07559_ (
  .A1(_02348_),
  .A2(_02349_),
  .ZN(_02350_)
);

NAND2_X1 _07560_ (
  .A1(_02350_),
  .A2(_02328_),
  .ZN(_02351_)
);

NAND2_X1 _07561_ (
  .A1(_02341_),
  .A2(\sresult[24][6] ),
  .ZN(_02352_)
);

NAND2_X1 _07562_ (
  .A1(_02351_),
  .A2(_02352_),
  .ZN(_00294_)
);

NAND2_X1 _07563_ (
  .A1(_02336_),
  .A2(\sresult[23][7] ),
  .ZN(_02353_)
);

NAND2_X1 _07564_ (
  .A1(_02325_),
  .A2(din_44[7]),
  .ZN(_02354_)
);

NAND2_X1 _07565_ (
  .A1(_02353_),
  .A2(_02354_),
  .ZN(_02355_)
);

NAND2_X1 _07566_ (
  .A1(_02355_),
  .A2(_02328_),
  .ZN(_02356_)
);

NAND2_X1 _07567_ (
  .A1(_02341_),
  .A2(\sresult[24][7] ),
  .ZN(_02357_)
);

NAND2_X1 _07568_ (
  .A1(_02356_),
  .A2(_02357_),
  .ZN(_00295_)
);

NAND2_X1 _07569_ (
  .A1(_02336_),
  .A2(\sresult[23][8] ),
  .ZN(_02358_)
);

NAND2_X1 _07570_ (
  .A1(_02325_),
  .A2(din_44[8]),
  .ZN(_02359_)
);

NAND2_X1 _07571_ (
  .A1(_02358_),
  .A2(_02359_),
  .ZN(_02360_)
);

NAND2_X1 _07572_ (
  .A1(_02360_),
  .A2(_02328_),
  .ZN(_02361_)
);

NAND2_X1 _07573_ (
  .A1(_02341_),
  .A2(\sresult[24][8] ),
  .ZN(_02362_)
);

NAND2_X1 _07574_ (
  .A1(_02361_),
  .A2(_02362_),
  .ZN(_00296_)
);

NAND2_X1 _07575_ (
  .A1(_02336_),
  .A2(\sresult[23][9] ),
  .ZN(_02363_)
);

NAND2_X1 _07576_ (
  .A1(_02325_),
  .A2(din_44[9]),
  .ZN(_02364_)
);

NAND2_X1 _07577_ (
  .A1(_02363_),
  .A2(_02364_),
  .ZN(_02365_)
);

NAND2_X1 _07578_ (
  .A1(_02365_),
  .A2(_02328_),
  .ZN(_02366_)
);

NAND2_X1 _07579_ (
  .A1(_02341_),
  .A2(\sresult[24][9] ),
  .ZN(_02367_)
);

NAND2_X1 _07580_ (
  .A1(_02366_),
  .A2(_02367_),
  .ZN(_00297_)
);

NAND2_X1 _07581_ (
  .A1(_02336_),
  .A2(\sresult[23][10] ),
  .ZN(_02368_)
);

NAND2_X1 _07582_ (
  .A1(_02325_),
  .A2(din_44[10]),
  .ZN(_02369_)
);

NAND2_X1 _07583_ (
  .A1(_02368_),
  .A2(_02369_),
  .ZN(_02370_)
);

NAND2_X1 _07584_ (
  .A1(_02370_),
  .A2(_02328_),
  .ZN(_02371_)
);

NAND2_X1 _07585_ (
  .A1(_02341_),
  .A2(\sresult[24][10] ),
  .ZN(_02372_)
);

NAND2_X1 _07586_ (
  .A1(_02371_),
  .A2(_02372_),
  .ZN(_00298_)
);

NAND2_X1 _07587_ (
  .A1(_02336_),
  .A2(\sresult[23][11] ),
  .ZN(_02373_)
);

NAND2_X1 _07588_ (
  .A1(_02325_),
  .A2(din_44[11]),
  .ZN(_02374_)
);

NAND2_X1 _07589_ (
  .A1(_02373_),
  .A2(_02374_),
  .ZN(_02375_)
);

NAND2_X1 _07590_ (
  .A1(_02375_),
  .A2(_02328_),
  .ZN(_02376_)
);

NAND2_X1 _07591_ (
  .A1(_02341_),
  .A2(\sresult[24][11] ),
  .ZN(_02377_)
);

NAND2_X1 _07592_ (
  .A1(_02376_),
  .A2(_02377_),
  .ZN(_00299_)
);

NAND2_X1 _07593_ (
  .A1(_02336_),
  .A2(\sresult[24][0] ),
  .ZN(_02378_)
);

BUF_X4 _07594_ (
  .A(_02107_),
  .Z(_02379_)
);

NAND2_X1 _07595_ (
  .A1(_02379_),
  .A2(din_53[0]),
  .ZN(_02380_)
);

NAND2_X1 _07596_ (
  .A1(_02378_),
  .A2(_02380_),
  .ZN(_02381_)
);

BUF_X2 _07597_ (
  .A(_02000_),
  .Z(_02382_)
);

NAND2_X1 _07598_ (
  .A1(_02381_),
  .A2(_02382_),
  .ZN(_02383_)
);

NAND2_X1 _07599_ (
  .A1(_02341_),
  .A2(\sresult[25][0] ),
  .ZN(_02384_)
);

NAND2_X1 _07600_ (
  .A1(_02383_),
  .A2(_02384_),
  .ZN(_00300_)
);

NAND2_X1 _07601_ (
  .A1(_02336_),
  .A2(\sresult[24][1] ),
  .ZN(_02385_)
);

NAND2_X1 _07602_ (
  .A1(_02379_),
  .A2(din_53[1]),
  .ZN(_02386_)
);

NAND2_X1 _07603_ (
  .A1(_02385_),
  .A2(_02386_),
  .ZN(_02387_)
);

NAND2_X1 _07604_ (
  .A1(_02387_),
  .A2(_02382_),
  .ZN(_02388_)
);

NAND2_X1 _07605_ (
  .A1(_02341_),
  .A2(\sresult[25][1] ),
  .ZN(_02389_)
);

NAND2_X1 _07606_ (
  .A1(_02388_),
  .A2(_02389_),
  .ZN(_00301_)
);

BUF_X4 _07607_ (
  .A(_02063_),
  .Z(_02390_)
);

NAND2_X1 _07608_ (
  .A1(_02390_),
  .A2(\sresult[24][2] ),
  .ZN(_02391_)
);

NAND2_X1 _07609_ (
  .A1(_02379_),
  .A2(din_53[2]),
  .ZN(_02392_)
);

NAND2_X1 _07610_ (
  .A1(_02391_),
  .A2(_02392_),
  .ZN(_02393_)
);

NAND2_X1 _07611_ (
  .A1(_02393_),
  .A2(_02382_),
  .ZN(_02394_)
);

BUF_X1 _07612_ (
  .A(_02124_),
  .Z(_02395_)
);

NAND2_X1 _07613_ (
  .A1(_02395_),
  .A2(\sresult[25][2] ),
  .ZN(_02396_)
);

NAND2_X1 _07614_ (
  .A1(_02394_),
  .A2(_02396_),
  .ZN(_00302_)
);

NAND2_X1 _07615_ (
  .A1(_02390_),
  .A2(\sresult[24][3] ),
  .ZN(_02397_)
);

NAND2_X1 _07616_ (
  .A1(_02379_),
  .A2(din_53[3]),
  .ZN(_02398_)
);

NAND2_X1 _07617_ (
  .A1(_02397_),
  .A2(_02398_),
  .ZN(_02399_)
);

NAND2_X1 _07618_ (
  .A1(_02399_),
  .A2(_02382_),
  .ZN(_02400_)
);

NAND2_X1 _07619_ (
  .A1(_02395_),
  .A2(\sresult[25][3] ),
  .ZN(_02401_)
);

NAND2_X1 _07620_ (
  .A1(_02400_),
  .A2(_02401_),
  .ZN(_00303_)
);

NAND2_X1 _07621_ (
  .A1(_02390_),
  .A2(\sresult[24][4] ),
  .ZN(_02402_)
);

NAND2_X1 _07622_ (
  .A1(_02379_),
  .A2(din_53[4]),
  .ZN(_02403_)
);

NAND2_X1 _07623_ (
  .A1(_02402_),
  .A2(_02403_),
  .ZN(_02404_)
);

NAND2_X1 _07624_ (
  .A1(_02404_),
  .A2(_02382_),
  .ZN(_02405_)
);

NAND2_X1 _07625_ (
  .A1(_02395_),
  .A2(\sresult[25][4] ),
  .ZN(_02406_)
);

NAND2_X1 _07626_ (
  .A1(_02405_),
  .A2(_02406_),
  .ZN(_00304_)
);

NAND2_X1 _07627_ (
  .A1(_02390_),
  .A2(\sresult[24][5] ),
  .ZN(_02407_)
);

NAND2_X1 _07628_ (
  .A1(_02379_),
  .A2(din_53[5]),
  .ZN(_02408_)
);

NAND2_X1 _07629_ (
  .A1(_02407_),
  .A2(_02408_),
  .ZN(_02409_)
);

NAND2_X1 _07630_ (
  .A1(_02409_),
  .A2(_02382_),
  .ZN(_02410_)
);

NAND2_X1 _07631_ (
  .A1(_02395_),
  .A2(\sresult[25][5] ),
  .ZN(_02411_)
);

NAND2_X1 _07632_ (
  .A1(_02410_),
  .A2(_02411_),
  .ZN(_00305_)
);

NAND2_X1 _07633_ (
  .A1(_02390_),
  .A2(\sresult[24][6] ),
  .ZN(_02412_)
);

NAND2_X1 _07634_ (
  .A1(_02379_),
  .A2(din_53[6]),
  .ZN(_02413_)
);

NAND2_X1 _07635_ (
  .A1(_02412_),
  .A2(_02413_),
  .ZN(_02414_)
);

NAND2_X1 _07636_ (
  .A1(_02414_),
  .A2(_02382_),
  .ZN(_02415_)
);

NAND2_X1 _07637_ (
  .A1(_02395_),
  .A2(\sresult[25][6] ),
  .ZN(_02416_)
);

NAND2_X1 _07638_ (
  .A1(_02415_),
  .A2(_02416_),
  .ZN(_00306_)
);

NAND2_X1 _07639_ (
  .A1(_02390_),
  .A2(\sresult[24][7] ),
  .ZN(_02417_)
);

NAND2_X1 _07640_ (
  .A1(_02379_),
  .A2(din_53[7]),
  .ZN(_02418_)
);

NAND2_X1 _07641_ (
  .A1(_02417_),
  .A2(_02418_),
  .ZN(_02419_)
);

NAND2_X1 _07642_ (
  .A1(_02419_),
  .A2(_02382_),
  .ZN(_02420_)
);

NAND2_X1 _07643_ (
  .A1(_02395_),
  .A2(\sresult[25][7] ),
  .ZN(_02421_)
);

NAND2_X1 _07644_ (
  .A1(_02420_),
  .A2(_02421_),
  .ZN(_00307_)
);

NAND2_X1 _07645_ (
  .A1(_02390_),
  .A2(\sresult[24][8] ),
  .ZN(_02422_)
);

NAND2_X1 _07646_ (
  .A1(_02379_),
  .A2(din_53[8]),
  .ZN(_02423_)
);

NAND2_X1 _07647_ (
  .A1(_02422_),
  .A2(_02423_),
  .ZN(_02424_)
);

NAND2_X1 _07648_ (
  .A1(_02424_),
  .A2(_02382_),
  .ZN(_02425_)
);

NAND2_X1 _07649_ (
  .A1(_02395_),
  .A2(\sresult[25][8] ),
  .ZN(_02426_)
);

NAND2_X1 _07650_ (
  .A1(_02425_),
  .A2(_02426_),
  .ZN(_00308_)
);

NAND2_X1 _07651_ (
  .A1(_02390_),
  .A2(\sresult[24][9] ),
  .ZN(_02427_)
);

NAND2_X1 _07652_ (
  .A1(_02379_),
  .A2(din_53[9]),
  .ZN(_02428_)
);

NAND2_X1 _07653_ (
  .A1(_02427_),
  .A2(_02428_),
  .ZN(_02429_)
);

NAND2_X1 _07654_ (
  .A1(_02429_),
  .A2(_02382_),
  .ZN(_02430_)
);

NAND2_X1 _07655_ (
  .A1(_02395_),
  .A2(\sresult[25][9] ),
  .ZN(_02431_)
);

NAND2_X1 _07656_ (
  .A1(_02430_),
  .A2(_02431_),
  .ZN(_00309_)
);

NAND2_X1 _07657_ (
  .A1(_02390_),
  .A2(\sresult[24][10] ),
  .ZN(_02432_)
);

BUF_X4 _07658_ (
  .A(_02107_),
  .Z(_02433_)
);

NAND2_X1 _07659_ (
  .A1(_02433_),
  .A2(din_53[10]),
  .ZN(_02434_)
);

NAND2_X1 _07660_ (
  .A1(_02432_),
  .A2(_02434_),
  .ZN(_02435_)
);

BUF_X2 _07661_ (
  .A(_02000_),
  .Z(_02436_)
);

NAND2_X1 _07662_ (
  .A1(_02435_),
  .A2(_02436_),
  .ZN(_02437_)
);

NAND2_X1 _07663_ (
  .A1(_02395_),
  .A2(\sresult[25][10] ),
  .ZN(_02438_)
);

NAND2_X1 _07664_ (
  .A1(_02437_),
  .A2(_02438_),
  .ZN(_00310_)
);

NAND2_X1 _07665_ (
  .A1(_02390_),
  .A2(\sresult[24][11] ),
  .ZN(_02439_)
);

NAND2_X1 _07666_ (
  .A1(_02433_),
  .A2(din_53[11]),
  .ZN(_02440_)
);

NAND2_X1 _07667_ (
  .A1(_02439_),
  .A2(_02440_),
  .ZN(_02441_)
);

NAND2_X1 _07668_ (
  .A1(_02441_),
  .A2(_02436_),
  .ZN(_02442_)
);

NAND2_X1 _07669_ (
  .A1(_02395_),
  .A2(\sresult[25][11] ),
  .ZN(_02443_)
);

NAND2_X1 _07670_ (
  .A1(_02442_),
  .A2(_02443_),
  .ZN(_00311_)
);

BUF_X4 _07671_ (
  .A(_02063_),
  .Z(_02444_)
);

NAND2_X1 _07672_ (
  .A1(_02444_),
  .A2(\sresult[25][0] ),
  .ZN(_02445_)
);

NAND2_X1 _07673_ (
  .A1(_02433_),
  .A2(din_62[0]),
  .ZN(_02446_)
);

NAND2_X1 _07674_ (
  .A1(_02445_),
  .A2(_02446_),
  .ZN(_02447_)
);

NAND2_X1 _07675_ (
  .A1(_02447_),
  .A2(_02436_),
  .ZN(_02448_)
);

BUF_X1 _07676_ (
  .A(_02124_),
  .Z(_02449_)
);

NAND2_X1 _07677_ (
  .A1(_02449_),
  .A2(\sresult[26][0] ),
  .ZN(_02450_)
);

NAND2_X1 _07678_ (
  .A1(_02448_),
  .A2(_02450_),
  .ZN(_00312_)
);

NAND2_X1 _07679_ (
  .A1(_02444_),
  .A2(\sresult[25][1] ),
  .ZN(_02451_)
);

NAND2_X1 _07680_ (
  .A1(_02433_),
  .A2(din_62[1]),
  .ZN(_02452_)
);

NAND2_X1 _07681_ (
  .A1(_02451_),
  .A2(_02452_),
  .ZN(_02453_)
);

NAND2_X1 _07682_ (
  .A1(_02453_),
  .A2(_02436_),
  .ZN(_02454_)
);

NAND2_X1 _07683_ (
  .A1(_02449_),
  .A2(\sresult[26][1] ),
  .ZN(_02455_)
);

NAND2_X1 _07684_ (
  .A1(_02454_),
  .A2(_02455_),
  .ZN(_00313_)
);

NAND2_X1 _07685_ (
  .A1(_02444_),
  .A2(\sresult[25][2] ),
  .ZN(_02456_)
);

NAND2_X1 _07686_ (
  .A1(_02433_),
  .A2(din_62[2]),
  .ZN(_02457_)
);

NAND2_X1 _07687_ (
  .A1(_02456_),
  .A2(_02457_),
  .ZN(_02458_)
);

NAND2_X1 _07688_ (
  .A1(_02458_),
  .A2(_02436_),
  .ZN(_02459_)
);

NAND2_X1 _07689_ (
  .A1(_02449_),
  .A2(\sresult[26][2] ),
  .ZN(_02460_)
);

NAND2_X1 _07690_ (
  .A1(_02459_),
  .A2(_02460_),
  .ZN(_00314_)
);

NAND2_X1 _07691_ (
  .A1(_02444_),
  .A2(\sresult[25][3] ),
  .ZN(_02461_)
);

NAND2_X1 _07692_ (
  .A1(_02433_),
  .A2(din_62[3]),
  .ZN(_02462_)
);

NAND2_X1 _07693_ (
  .A1(_02461_),
  .A2(_02462_),
  .ZN(_02463_)
);

NAND2_X1 _07694_ (
  .A1(_02463_),
  .A2(_02436_),
  .ZN(_02464_)
);

NAND2_X1 _07695_ (
  .A1(_02449_),
  .A2(\sresult[26][3] ),
  .ZN(_02465_)
);

NAND2_X1 _07696_ (
  .A1(_02464_),
  .A2(_02465_),
  .ZN(_00315_)
);

NAND2_X1 _07697_ (
  .A1(_02444_),
  .A2(\sresult[25][4] ),
  .ZN(_02466_)
);

NAND2_X1 _07698_ (
  .A1(_02433_),
  .A2(din_62[4]),
  .ZN(_02467_)
);

NAND2_X1 _07699_ (
  .A1(_02466_),
  .A2(_02467_),
  .ZN(_02468_)
);

NAND2_X1 _07700_ (
  .A1(_02468_),
  .A2(_02436_),
  .ZN(_02469_)
);

NAND2_X1 _07701_ (
  .A1(_02449_),
  .A2(\sresult[26][4] ),
  .ZN(_02470_)
);

NAND2_X1 _07702_ (
  .A1(_02469_),
  .A2(_02470_),
  .ZN(_00316_)
);

NAND2_X1 _07703_ (
  .A1(_02444_),
  .A2(\sresult[25][5] ),
  .ZN(_02471_)
);

NAND2_X1 _07704_ (
  .A1(_02433_),
  .A2(din_62[5]),
  .ZN(_02472_)
);

NAND2_X1 _07705_ (
  .A1(_02471_),
  .A2(_02472_),
  .ZN(_02473_)
);

NAND2_X1 _07706_ (
  .A1(_02473_),
  .A2(_02436_),
  .ZN(_02474_)
);

NAND2_X1 _07707_ (
  .A1(_02449_),
  .A2(\sresult[26][5] ),
  .ZN(_02475_)
);

NAND2_X1 _07708_ (
  .A1(_02474_),
  .A2(_02475_),
  .ZN(_00317_)
);

NAND2_X1 _07709_ (
  .A1(_02444_),
  .A2(\sresult[25][6] ),
  .ZN(_02476_)
);

NAND2_X1 _07710_ (
  .A1(_02433_),
  .A2(din_62[6]),
  .ZN(_02477_)
);

NAND2_X1 _07711_ (
  .A1(_02476_),
  .A2(_02477_),
  .ZN(_02478_)
);

NAND2_X1 _07712_ (
  .A1(_02478_),
  .A2(_02436_),
  .ZN(_02479_)
);

NAND2_X1 _07713_ (
  .A1(_02449_),
  .A2(\sresult[26][6] ),
  .ZN(_02480_)
);

NAND2_X1 _07714_ (
  .A1(_02479_),
  .A2(_02480_),
  .ZN(_00318_)
);

NAND2_X1 _07715_ (
  .A1(_02444_),
  .A2(\sresult[25][7] ),
  .ZN(_02481_)
);

NAND2_X1 _07716_ (
  .A1(_02433_),
  .A2(din_62[7]),
  .ZN(_02482_)
);

NAND2_X1 _07717_ (
  .A1(_02481_),
  .A2(_02482_),
  .ZN(_02483_)
);

NAND2_X1 _07718_ (
  .A1(_02483_),
  .A2(_02436_),
  .ZN(_02484_)
);

NAND2_X1 _07719_ (
  .A1(_02449_),
  .A2(\sresult[26][7] ),
  .ZN(_02485_)
);

NAND2_X1 _07720_ (
  .A1(_02484_),
  .A2(_02485_),
  .ZN(_00319_)
);

NAND2_X1 _07721_ (
  .A1(_02444_),
  .A2(\sresult[25][8] ),
  .ZN(_02486_)
);

BUF_X4 _07722_ (
  .A(_02107_),
  .Z(_02487_)
);

NAND2_X1 _07723_ (
  .A1(_02487_),
  .A2(din_62[8]),
  .ZN(_02488_)
);

NAND2_X1 _07724_ (
  .A1(_02486_),
  .A2(_02488_),
  .ZN(_02489_)
);

BUF_X2 _07725_ (
  .A(_02000_),
  .Z(_02490_)
);

NAND2_X1 _07726_ (
  .A1(_02489_),
  .A2(_02490_),
  .ZN(_02491_)
);

NAND2_X1 _07727_ (
  .A1(_02449_),
  .A2(\sresult[26][8] ),
  .ZN(_02492_)
);

NAND2_X1 _07728_ (
  .A1(_02491_),
  .A2(_02492_),
  .ZN(_00320_)
);

NAND2_X1 _07729_ (
  .A1(_02444_),
  .A2(\sresult[25][9] ),
  .ZN(_02493_)
);

NAND2_X1 _07730_ (
  .A1(_02487_),
  .A2(din_62[9]),
  .ZN(_02494_)
);

NAND2_X1 _07731_ (
  .A1(_02493_),
  .A2(_02494_),
  .ZN(_02495_)
);

NAND2_X1 _07732_ (
  .A1(_02495_),
  .A2(_02490_),
  .ZN(_02496_)
);

NAND2_X1 _07733_ (
  .A1(_02449_),
  .A2(\sresult[26][9] ),
  .ZN(_02497_)
);

NAND2_X1 _07734_ (
  .A1(_02496_),
  .A2(_02497_),
  .ZN(_00321_)
);

BUF_X4 _07735_ (
  .A(_02063_),
  .Z(_02498_)
);

NAND2_X1 _07736_ (
  .A1(_02498_),
  .A2(\sresult[25][10] ),
  .ZN(_02499_)
);

NAND2_X1 _07737_ (
  .A1(_02487_),
  .A2(din_62[10]),
  .ZN(_02500_)
);

NAND2_X1 _07738_ (
  .A1(_02499_),
  .A2(_02500_),
  .ZN(_02501_)
);

NAND2_X1 _07739_ (
  .A1(_02501_),
  .A2(_02490_),
  .ZN(_02502_)
);

BUF_X1 _07740_ (
  .A(_02124_),
  .Z(_02503_)
);

NAND2_X1 _07741_ (
  .A1(_02503_),
  .A2(\sresult[26][10] ),
  .ZN(_02504_)
);

NAND2_X1 _07742_ (
  .A1(_02502_),
  .A2(_02504_),
  .ZN(_00322_)
);

NAND2_X1 _07743_ (
  .A1(_02498_),
  .A2(\sresult[25][11] ),
  .ZN(_02505_)
);

NAND2_X1 _07744_ (
  .A1(_02487_),
  .A2(din_62[11]),
  .ZN(_02506_)
);

NAND2_X1 _07745_ (
  .A1(_02505_),
  .A2(_02506_),
  .ZN(_02507_)
);

NAND2_X1 _07746_ (
  .A1(_02507_),
  .A2(_02490_),
  .ZN(_02508_)
);

NAND2_X1 _07747_ (
  .A1(_02503_),
  .A2(\sresult[26][11] ),
  .ZN(_02509_)
);

NAND2_X1 _07748_ (
  .A1(_02508_),
  .A2(_02509_),
  .ZN(_00323_)
);

NAND2_X1 _07749_ (
  .A1(_02498_),
  .A2(\sresult[26][0] ),
  .ZN(_02510_)
);

NAND2_X1 _07750_ (
  .A1(_02487_),
  .A2(din_71[0]),
  .ZN(_02511_)
);

NAND2_X1 _07751_ (
  .A1(_02510_),
  .A2(_02511_),
  .ZN(_02512_)
);

NAND2_X1 _07752_ (
  .A1(_02512_),
  .A2(_02490_),
  .ZN(_02513_)
);

NAND2_X1 _07753_ (
  .A1(_02503_),
  .A2(\sresult[27][0] ),
  .ZN(_02514_)
);

NAND2_X1 _07754_ (
  .A1(_02513_),
  .A2(_02514_),
  .ZN(_00324_)
);

NAND2_X1 _07755_ (
  .A1(_02498_),
  .A2(\sresult[26][1] ),
  .ZN(_02515_)
);

NAND2_X1 _07756_ (
  .A1(_02487_),
  .A2(din_71[1]),
  .ZN(_02516_)
);

NAND2_X1 _07757_ (
  .A1(_02515_),
  .A2(_02516_),
  .ZN(_02517_)
);

NAND2_X1 _07758_ (
  .A1(_02517_),
  .A2(_02490_),
  .ZN(_02518_)
);

NAND2_X1 _07759_ (
  .A1(_02503_),
  .A2(\sresult[27][1] ),
  .ZN(_02519_)
);

NAND2_X1 _07760_ (
  .A1(_02518_),
  .A2(_02519_),
  .ZN(_00325_)
);

NAND2_X1 _07761_ (
  .A1(_02498_),
  .A2(\sresult[26][2] ),
  .ZN(_02520_)
);

NAND2_X1 _07762_ (
  .A1(_02487_),
  .A2(din_71[2]),
  .ZN(_02521_)
);

NAND2_X1 _07763_ (
  .A1(_02520_),
  .A2(_02521_),
  .ZN(_02522_)
);

NAND2_X1 _07764_ (
  .A1(_02522_),
  .A2(_02490_),
  .ZN(_02523_)
);

NAND2_X1 _07765_ (
  .A1(_02503_),
  .A2(\sresult[27][2] ),
  .ZN(_02524_)
);

NAND2_X1 _07766_ (
  .A1(_02523_),
  .A2(_02524_),
  .ZN(_00326_)
);

NAND2_X1 _07767_ (
  .A1(_02498_),
  .A2(\sresult[26][3] ),
  .ZN(_02525_)
);

NAND2_X1 _07768_ (
  .A1(_02487_),
  .A2(din_71[3]),
  .ZN(_02526_)
);

NAND2_X1 _07769_ (
  .A1(_02525_),
  .A2(_02526_),
  .ZN(_02527_)
);

NAND2_X1 _07770_ (
  .A1(_02527_),
  .A2(_02490_),
  .ZN(_02528_)
);

NAND2_X1 _07771_ (
  .A1(_02503_),
  .A2(\sresult[27][3] ),
  .ZN(_02529_)
);

NAND2_X1 _07772_ (
  .A1(_02528_),
  .A2(_02529_),
  .ZN(_00327_)
);

NAND2_X1 _07773_ (
  .A1(_02498_),
  .A2(\sresult[26][4] ),
  .ZN(_02530_)
);

NAND2_X1 _07774_ (
  .A1(_02487_),
  .A2(din_71[4]),
  .ZN(_02531_)
);

NAND2_X1 _07775_ (
  .A1(_02530_),
  .A2(_02531_),
  .ZN(_02532_)
);

NAND2_X1 _07776_ (
  .A1(_02532_),
  .A2(_02490_),
  .ZN(_02533_)
);

NAND2_X1 _07777_ (
  .A1(_02503_),
  .A2(\sresult[27][4] ),
  .ZN(_02534_)
);

NAND2_X1 _07778_ (
  .A1(_02533_),
  .A2(_02534_),
  .ZN(_00328_)
);

NAND2_X1 _07779_ (
  .A1(_02498_),
  .A2(\sresult[26][5] ),
  .ZN(_02535_)
);

NAND2_X1 _07780_ (
  .A1(_02487_),
  .A2(din_71[5]),
  .ZN(_02536_)
);

NAND2_X1 _07781_ (
  .A1(_02535_),
  .A2(_02536_),
  .ZN(_02537_)
);

NAND2_X1 _07782_ (
  .A1(_02537_),
  .A2(_02490_),
  .ZN(_02538_)
);

NAND2_X1 _07783_ (
  .A1(_02503_),
  .A2(\sresult[27][5] ),
  .ZN(_02539_)
);

NAND2_X1 _07784_ (
  .A1(_02538_),
  .A2(_02539_),
  .ZN(_00329_)
);

NAND2_X1 _07785_ (
  .A1(_02498_),
  .A2(\sresult[26][6] ),
  .ZN(_02540_)
);

BUF_X4 _07786_ (
  .A(_02107_),
  .Z(_02541_)
);

NAND2_X1 _07787_ (
  .A1(_02541_),
  .A2(din_71[6]),
  .ZN(_02542_)
);

NAND2_X1 _07788_ (
  .A1(_02540_),
  .A2(_02542_),
  .ZN(_02543_)
);

BUF_X4 _07789_ (
  .A(_00911_),
  .Z(_02544_)
);

BUF_X2 _07790_ (
  .A(_02544_),
  .Z(_02545_)
);

NAND2_X1 _07791_ (
  .A1(_02543_),
  .A2(_02545_),
  .ZN(_02546_)
);

NAND2_X1 _07792_ (
  .A1(_02503_),
  .A2(\sresult[27][6] ),
  .ZN(_02547_)
);

NAND2_X1 _07793_ (
  .A1(_02546_),
  .A2(_02547_),
  .ZN(_00330_)
);

NAND2_X1 _07794_ (
  .A1(_02498_),
  .A2(\sresult[26][7] ),
  .ZN(_02548_)
);

NAND2_X1 _07795_ (
  .A1(_02541_),
  .A2(din_71[7]),
  .ZN(_02549_)
);

NAND2_X1 _07796_ (
  .A1(_02548_),
  .A2(_02549_),
  .ZN(_02550_)
);

NAND2_X1 _07797_ (
  .A1(_02550_),
  .A2(_02545_),
  .ZN(_02551_)
);

NAND2_X1 _07798_ (
  .A1(_02503_),
  .A2(\sresult[27][7] ),
  .ZN(_02552_)
);

NAND2_X1 _07799_ (
  .A1(_02551_),
  .A2(_02552_),
  .ZN(_00331_)
);

BUF_X4 _07800_ (
  .A(_02063_),
  .Z(_02553_)
);

NAND2_X1 _07801_ (
  .A1(_02553_),
  .A2(\sresult[26][8] ),
  .ZN(_02554_)
);

NAND2_X1 _07802_ (
  .A1(_02541_),
  .A2(din_71[8]),
  .ZN(_02555_)
);

NAND2_X1 _07803_ (
  .A1(_02554_),
  .A2(_02555_),
  .ZN(_02556_)
);

NAND2_X1 _07804_ (
  .A1(_02556_),
  .A2(_02545_),
  .ZN(_02557_)
);

BUF_X1 _07805_ (
  .A(_02124_),
  .Z(_02558_)
);

NAND2_X1 _07806_ (
  .A1(_02558_),
  .A2(\sresult[27][8] ),
  .ZN(_02559_)
);

NAND2_X1 _07807_ (
  .A1(_02557_),
  .A2(_02559_),
  .ZN(_00332_)
);

NAND2_X1 _07808_ (
  .A1(_02553_),
  .A2(\sresult[26][9] ),
  .ZN(_02560_)
);

NAND2_X1 _07809_ (
  .A1(_02541_),
  .A2(din_71[9]),
  .ZN(_02561_)
);

NAND2_X1 _07810_ (
  .A1(_02560_),
  .A2(_02561_),
  .ZN(_02562_)
);

NAND2_X1 _07811_ (
  .A1(_02562_),
  .A2(_02545_),
  .ZN(_02563_)
);

NAND2_X1 _07812_ (
  .A1(_02558_),
  .A2(\sresult[27][9] ),
  .ZN(_02564_)
);

NAND2_X1 _07813_ (
  .A1(_02563_),
  .A2(_02564_),
  .ZN(_00333_)
);

NAND2_X1 _07814_ (
  .A1(_02553_),
  .A2(\sresult[26][10] ),
  .ZN(_02565_)
);

NAND2_X1 _07815_ (
  .A1(_02541_),
  .A2(din_71[10]),
  .ZN(_02566_)
);

NAND2_X1 _07816_ (
  .A1(_02565_),
  .A2(_02566_),
  .ZN(_02567_)
);

NAND2_X1 _07817_ (
  .A1(_02567_),
  .A2(_02545_),
  .ZN(_02568_)
);

NAND2_X1 _07818_ (
  .A1(_02558_),
  .A2(\sresult[27][10] ),
  .ZN(_02569_)
);

NAND2_X1 _07819_ (
  .A1(_02568_),
  .A2(_02569_),
  .ZN(_00334_)
);

NAND2_X1 _07820_ (
  .A1(_02553_),
  .A2(\sresult[26][11] ),
  .ZN(_02570_)
);

NAND2_X1 _07821_ (
  .A1(_02541_),
  .A2(din_71[11]),
  .ZN(_02571_)
);

NAND2_X1 _07822_ (
  .A1(_02570_),
  .A2(_02571_),
  .ZN(_02572_)
);

NAND2_X1 _07823_ (
  .A1(_02572_),
  .A2(_02545_),
  .ZN(_02573_)
);

NAND2_X1 _07824_ (
  .A1(_02558_),
  .A2(\sresult[27][11] ),
  .ZN(_02574_)
);

NAND2_X1 _07825_ (
  .A1(_02573_),
  .A2(_02574_),
  .ZN(_00335_)
);

NAND2_X1 _07826_ (
  .A1(_02553_),
  .A2(\sresult[27][0] ),
  .ZN(_02575_)
);

NAND2_X1 _07827_ (
  .A1(_02541_),
  .A2(din_70[0]),
  .ZN(_02576_)
);

NAND2_X1 _07828_ (
  .A1(_02575_),
  .A2(_02576_),
  .ZN(_02577_)
);

NAND2_X1 _07829_ (
  .A1(_02577_),
  .A2(_02545_),
  .ZN(_02578_)
);

NAND2_X1 _07830_ (
  .A1(_02558_),
  .A2(\sresult[28][0] ),
  .ZN(_02579_)
);

NAND2_X1 _07831_ (
  .A1(_02578_),
  .A2(_02579_),
  .ZN(_00336_)
);

NAND2_X1 _07832_ (
  .A1(_02553_),
  .A2(\sresult[27][1] ),
  .ZN(_02580_)
);

NAND2_X1 _07833_ (
  .A1(_02541_),
  .A2(din_70[1]),
  .ZN(_02581_)
);

NAND2_X1 _07834_ (
  .A1(_02580_),
  .A2(_02581_),
  .ZN(_02582_)
);

NAND2_X1 _07835_ (
  .A1(_02582_),
  .A2(_02545_),
  .ZN(_02583_)
);

NAND2_X1 _07836_ (
  .A1(_02558_),
  .A2(\sresult[28][1] ),
  .ZN(_02584_)
);

NAND2_X1 _07837_ (
  .A1(_02583_),
  .A2(_02584_),
  .ZN(_00337_)
);

NAND2_X1 _07838_ (
  .A1(_02553_),
  .A2(\sresult[27][2] ),
  .ZN(_02585_)
);

NAND2_X1 _07839_ (
  .A1(_02541_),
  .A2(din_70[2]),
  .ZN(_02586_)
);

NAND2_X1 _07840_ (
  .A1(_02585_),
  .A2(_02586_),
  .ZN(_02587_)
);

NAND2_X1 _07841_ (
  .A1(_02587_),
  .A2(_02545_),
  .ZN(_02588_)
);

NAND2_X1 _07842_ (
  .A1(_02558_),
  .A2(\sresult[28][2] ),
  .ZN(_02589_)
);

NAND2_X1 _07843_ (
  .A1(_02588_),
  .A2(_02589_),
  .ZN(_00338_)
);

NAND2_X1 _07844_ (
  .A1(_02553_),
  .A2(\sresult[27][3] ),
  .ZN(_02590_)
);

NAND2_X1 _07845_ (
  .A1(_02541_),
  .A2(din_70[3]),
  .ZN(_02591_)
);

NAND2_X1 _07846_ (
  .A1(_02590_),
  .A2(_02591_),
  .ZN(_02592_)
);

NAND2_X1 _07847_ (
  .A1(_02592_),
  .A2(_02545_),
  .ZN(_02593_)
);

NAND2_X1 _07848_ (
  .A1(_02558_),
  .A2(\sresult[28][3] ),
  .ZN(_02594_)
);

NAND2_X1 _07849_ (
  .A1(_02593_),
  .A2(_02594_),
  .ZN(_00339_)
);

NAND2_X1 _07850_ (
  .A1(_02553_),
  .A2(\sresult[27][4] ),
  .ZN(_02595_)
);

BUF_X4 _07851_ (
  .A(_02107_),
  .Z(_02596_)
);

NAND2_X1 _07852_ (
  .A1(_02596_),
  .A2(din_70[4]),
  .ZN(_02597_)
);

NAND2_X1 _07853_ (
  .A1(_02595_),
  .A2(_02597_),
  .ZN(_02598_)
);

BUF_X2 _07854_ (
  .A(_02544_),
  .Z(_02599_)
);

NAND2_X1 _07855_ (
  .A1(_02598_),
  .A2(_02599_),
  .ZN(_02600_)
);

NAND2_X1 _07856_ (
  .A1(_02558_),
  .A2(\sresult[28][4] ),
  .ZN(_02601_)
);

NAND2_X1 _07857_ (
  .A1(_02600_),
  .A2(_02601_),
  .ZN(_00340_)
);

NAND2_X1 _07858_ (
  .A1(_02553_),
  .A2(\sresult[27][5] ),
  .ZN(_02602_)
);

NAND2_X1 _07859_ (
  .A1(_02596_),
  .A2(din_70[5]),
  .ZN(_02603_)
);

NAND2_X1 _07860_ (
  .A1(_02602_),
  .A2(_02603_),
  .ZN(_02604_)
);

NAND2_X1 _07861_ (
  .A1(_02604_),
  .A2(_02599_),
  .ZN(_02605_)
);

NAND2_X1 _07862_ (
  .A1(_02558_),
  .A2(\sresult[28][5] ),
  .ZN(_02606_)
);

NAND2_X1 _07863_ (
  .A1(_02605_),
  .A2(_02606_),
  .ZN(_00341_)
);

BUF_X4 _07864_ (
  .A(_00800_),
  .Z(_02607_)
);

NAND2_X1 _07865_ (
  .A1(_02607_),
  .A2(\sresult[27][6] ),
  .ZN(_02608_)
);

NAND2_X1 _07866_ (
  .A1(_02596_),
  .A2(din_70[6]),
  .ZN(_02609_)
);

NAND2_X1 _07867_ (
  .A1(_02608_),
  .A2(_02609_),
  .ZN(_02610_)
);

NAND2_X1 _07868_ (
  .A1(_02610_),
  .A2(_02599_),
  .ZN(_02611_)
);

BUF_X1 _07869_ (
  .A(_02124_),
  .Z(_02612_)
);

NAND2_X1 _07870_ (
  .A1(_02612_),
  .A2(\sresult[28][6] ),
  .ZN(_02613_)
);

NAND2_X1 _07871_ (
  .A1(_02611_),
  .A2(_02613_),
  .ZN(_00342_)
);

NAND2_X1 _07872_ (
  .A1(_02607_),
  .A2(\sresult[27][7] ),
  .ZN(_02614_)
);

NAND2_X1 _07873_ (
  .A1(_02596_),
  .A2(din_70[7]),
  .ZN(_02615_)
);

NAND2_X1 _07874_ (
  .A1(_02614_),
  .A2(_02615_),
  .ZN(_02616_)
);

NAND2_X1 _07875_ (
  .A1(_02616_),
  .A2(_02599_),
  .ZN(_02617_)
);

NAND2_X1 _07876_ (
  .A1(_02612_),
  .A2(\sresult[28][7] ),
  .ZN(_02618_)
);

NAND2_X1 _07877_ (
  .A1(_02617_),
  .A2(_02618_),
  .ZN(_00343_)
);

NAND2_X1 _07878_ (
  .A1(_02607_),
  .A2(\sresult[27][8] ),
  .ZN(_02619_)
);

NAND2_X1 _07879_ (
  .A1(_02596_),
  .A2(din_70[8]),
  .ZN(_02620_)
);

NAND2_X1 _07880_ (
  .A1(_02619_),
  .A2(_02620_),
  .ZN(_02621_)
);

NAND2_X1 _07881_ (
  .A1(_02621_),
  .A2(_02599_),
  .ZN(_02622_)
);

NAND2_X1 _07882_ (
  .A1(_02612_),
  .A2(\sresult[28][8] ),
  .ZN(_02623_)
);

NAND2_X1 _07883_ (
  .A1(_02622_),
  .A2(_02623_),
  .ZN(_00344_)
);

NAND2_X1 _07884_ (
  .A1(_02607_),
  .A2(\sresult[27][9] ),
  .ZN(_02624_)
);

NAND2_X1 _07885_ (
  .A1(_02596_),
  .A2(din_70[9]),
  .ZN(_02625_)
);

NAND2_X1 _07886_ (
  .A1(_02624_),
  .A2(_02625_),
  .ZN(_02626_)
);

NAND2_X1 _07887_ (
  .A1(_02626_),
  .A2(_02599_),
  .ZN(_02627_)
);

NAND2_X1 _07888_ (
  .A1(_02612_),
  .A2(\sresult[28][9] ),
  .ZN(_02628_)
);

NAND2_X1 _07889_ (
  .A1(_02627_),
  .A2(_02628_),
  .ZN(_00345_)
);

NAND2_X1 _07890_ (
  .A1(_02607_),
  .A2(\sresult[27][10] ),
  .ZN(_02629_)
);

NAND2_X1 _07891_ (
  .A1(_02596_),
  .A2(din_70[10]),
  .ZN(_02630_)
);

NAND2_X1 _07892_ (
  .A1(_02629_),
  .A2(_02630_),
  .ZN(_02631_)
);

NAND2_X1 _07893_ (
  .A1(_02631_),
  .A2(_02599_),
  .ZN(_02632_)
);

NAND2_X1 _07894_ (
  .A1(_02612_),
  .A2(\sresult[28][10] ),
  .ZN(_02633_)
);

NAND2_X1 _07895_ (
  .A1(_02632_),
  .A2(_02633_),
  .ZN(_00346_)
);

NAND2_X1 _07896_ (
  .A1(_02607_),
  .A2(\sresult[27][11] ),
  .ZN(_02634_)
);

NAND2_X1 _07897_ (
  .A1(_02596_),
  .A2(din_70[11]),
  .ZN(_02635_)
);

NAND2_X1 _07898_ (
  .A1(_02634_),
  .A2(_02635_),
  .ZN(_02636_)
);

NAND2_X1 _07899_ (
  .A1(_02636_),
  .A2(_02599_),
  .ZN(_02637_)
);

NAND2_X1 _07900_ (
  .A1(_02612_),
  .A2(\sresult[28][11] ),
  .ZN(_02638_)
);

NAND2_X1 _07901_ (
  .A1(_02637_),
  .A2(_02638_),
  .ZN(_00347_)
);

NAND2_X1 _07902_ (
  .A1(_02607_),
  .A2(\sresult[28][0] ),
  .ZN(_02639_)
);

NAND2_X1 _07903_ (
  .A1(_02596_),
  .A2(din_61[0]),
  .ZN(_02640_)
);

NAND2_X1 _07904_ (
  .A1(_02639_),
  .A2(_02640_),
  .ZN(_02641_)
);

NAND2_X1 _07905_ (
  .A1(_02641_),
  .A2(_02599_),
  .ZN(_02642_)
);

NAND2_X1 _07906_ (
  .A1(_02612_),
  .A2(\sresult[29][0] ),
  .ZN(_02643_)
);

NAND2_X1 _07907_ (
  .A1(_02642_),
  .A2(_02643_),
  .ZN(_00348_)
);

NAND2_X1 _07908_ (
  .A1(_02607_),
  .A2(\sresult[28][1] ),
  .ZN(_02644_)
);

NAND2_X1 _07909_ (
  .A1(_02596_),
  .A2(din_61[1]),
  .ZN(_02645_)
);

NAND2_X1 _07910_ (
  .A1(_02644_),
  .A2(_02645_),
  .ZN(_02646_)
);

NAND2_X1 _07911_ (
  .A1(_02646_),
  .A2(_02599_),
  .ZN(_02647_)
);

NAND2_X1 _07912_ (
  .A1(_02612_),
  .A2(\sresult[29][1] ),
  .ZN(_02648_)
);

NAND2_X1 _07913_ (
  .A1(_02647_),
  .A2(_02648_),
  .ZN(_00349_)
);

NAND2_X1 _07914_ (
  .A1(_02607_),
  .A2(\sresult[28][2] ),
  .ZN(_02649_)
);

BUF_X8 _07915_ (
  .A(_00770_),
  .Z(_02650_)
);

BUF_X4 _07916_ (
  .A(_02650_),
  .Z(_02651_)
);

NAND2_X1 _07917_ (
  .A1(_02651_),
  .A2(din_61[2]),
  .ZN(_02652_)
);

NAND2_X1 _07918_ (
  .A1(_02649_),
  .A2(_02652_),
  .ZN(_02653_)
);

BUF_X2 _07919_ (
  .A(_02544_),
  .Z(_02654_)
);

NAND2_X1 _07920_ (
  .A1(_02653_),
  .A2(_02654_),
  .ZN(_02655_)
);

NAND2_X1 _07921_ (
  .A1(_02612_),
  .A2(\sresult[29][2] ),
  .ZN(_02656_)
);

NAND2_X1 _07922_ (
  .A1(_02655_),
  .A2(_02656_),
  .ZN(_00350_)
);

NAND2_X1 _07923_ (
  .A1(_02607_),
  .A2(\sresult[28][3] ),
  .ZN(_02657_)
);

NAND2_X1 _07924_ (
  .A1(_02651_),
  .A2(din_61[3]),
  .ZN(_02658_)
);

NAND2_X1 _07925_ (
  .A1(_02657_),
  .A2(_02658_),
  .ZN(_02659_)
);

NAND2_X1 _07926_ (
  .A1(_02659_),
  .A2(_02654_),
  .ZN(_02660_)
);

NAND2_X1 _07927_ (
  .A1(_02612_),
  .A2(\sresult[29][3] ),
  .ZN(_02661_)
);

NAND2_X1 _07928_ (
  .A1(_02660_),
  .A2(_02661_),
  .ZN(_00351_)
);

BUF_X4 _07929_ (
  .A(_00800_),
  .Z(_02662_)
);

NAND2_X1 _07930_ (
  .A1(_02662_),
  .A2(\sresult[28][4] ),
  .ZN(_02663_)
);

NAND2_X1 _07931_ (
  .A1(_02651_),
  .A2(din_61[4]),
  .ZN(_02664_)
);

NAND2_X1 _07932_ (
  .A1(_02663_),
  .A2(_02664_),
  .ZN(_02665_)
);

NAND2_X1 _07933_ (
  .A1(_02665_),
  .A2(_02654_),
  .ZN(_02666_)
);

BUF_X1 _07934_ (
  .A(_00811_),
  .Z(_02667_)
);

NAND2_X1 _07935_ (
  .A1(_02667_),
  .A2(\sresult[29][4] ),
  .ZN(_02668_)
);

NAND2_X1 _07936_ (
  .A1(_02666_),
  .A2(_02668_),
  .ZN(_00352_)
);

NAND2_X1 _07937_ (
  .A1(_02662_),
  .A2(\sresult[28][5] ),
  .ZN(_02669_)
);

NAND2_X1 _07938_ (
  .A1(_02651_),
  .A2(din_61[5]),
  .ZN(_02670_)
);

NAND2_X1 _07939_ (
  .A1(_02669_),
  .A2(_02670_),
  .ZN(_02671_)
);

NAND2_X1 _07940_ (
  .A1(_02671_),
  .A2(_02654_),
  .ZN(_02672_)
);

NAND2_X1 _07941_ (
  .A1(_02667_),
  .A2(\sresult[29][5] ),
  .ZN(_02673_)
);

NAND2_X1 _07942_ (
  .A1(_02672_),
  .A2(_02673_),
  .ZN(_00353_)
);

NAND2_X1 _07943_ (
  .A1(_02662_),
  .A2(\sresult[28][6] ),
  .ZN(_02674_)
);

NAND2_X1 _07944_ (
  .A1(_02651_),
  .A2(din_61[6]),
  .ZN(_02675_)
);

NAND2_X1 _07945_ (
  .A1(_02674_),
  .A2(_02675_),
  .ZN(_02676_)
);

NAND2_X1 _07946_ (
  .A1(_02676_),
  .A2(_02654_),
  .ZN(_02677_)
);

NAND2_X1 _07947_ (
  .A1(_02667_),
  .A2(\sresult[29][6] ),
  .ZN(_02678_)
);

NAND2_X1 _07948_ (
  .A1(_02677_),
  .A2(_02678_),
  .ZN(_00354_)
);

NAND2_X1 _07949_ (
  .A1(_02662_),
  .A2(\sresult[28][7] ),
  .ZN(_02679_)
);

NAND2_X1 _07950_ (
  .A1(_02651_),
  .A2(din_61[7]),
  .ZN(_02680_)
);

NAND2_X1 _07951_ (
  .A1(_02679_),
  .A2(_02680_),
  .ZN(_02681_)
);

NAND2_X1 _07952_ (
  .A1(_02681_),
  .A2(_02654_),
  .ZN(_02682_)
);

NAND2_X1 _07953_ (
  .A1(_02667_),
  .A2(\sresult[29][7] ),
  .ZN(_02683_)
);

NAND2_X1 _07954_ (
  .A1(_02682_),
  .A2(_02683_),
  .ZN(_00355_)
);

NAND2_X1 _07955_ (
  .A1(_02662_),
  .A2(\sresult[28][8] ),
  .ZN(_02684_)
);

NAND2_X1 _07956_ (
  .A1(_02651_),
  .A2(din_61[8]),
  .ZN(_02685_)
);

NAND2_X1 _07957_ (
  .A1(_02684_),
  .A2(_02685_),
  .ZN(_02686_)
);

NAND2_X1 _07958_ (
  .A1(_02686_),
  .A2(_02654_),
  .ZN(_02687_)
);

NAND2_X1 _07959_ (
  .A1(_02667_),
  .A2(\sresult[29][8] ),
  .ZN(_02688_)
);

NAND2_X1 _07960_ (
  .A1(_02687_),
  .A2(_02688_),
  .ZN(_00356_)
);

NAND2_X1 _07961_ (
  .A1(_02662_),
  .A2(\sresult[28][9] ),
  .ZN(_02689_)
);

NAND2_X1 _07962_ (
  .A1(_02651_),
  .A2(din_61[9]),
  .ZN(_02690_)
);

NAND2_X1 _07963_ (
  .A1(_02689_),
  .A2(_02690_),
  .ZN(_02691_)
);

NAND2_X1 _07964_ (
  .A1(_02691_),
  .A2(_02654_),
  .ZN(_02692_)
);

NAND2_X1 _07965_ (
  .A1(_02667_),
  .A2(\sresult[29][9] ),
  .ZN(_02693_)
);

NAND2_X1 _07966_ (
  .A1(_02692_),
  .A2(_02693_),
  .ZN(_00357_)
);

NAND2_X1 _07967_ (
  .A1(_02662_),
  .A2(\sresult[28][10] ),
  .ZN(_02694_)
);

NAND2_X1 _07968_ (
  .A1(_02651_),
  .A2(din_61[10]),
  .ZN(_02695_)
);

NAND2_X1 _07969_ (
  .A1(_02694_),
  .A2(_02695_),
  .ZN(_02696_)
);

NAND2_X1 _07970_ (
  .A1(_02696_),
  .A2(_02654_),
  .ZN(_02697_)
);

NAND2_X1 _07971_ (
  .A1(_02667_),
  .A2(\sresult[29][10] ),
  .ZN(_02698_)
);

NAND2_X1 _07972_ (
  .A1(_02697_),
  .A2(_02698_),
  .ZN(_00358_)
);

NAND2_X1 _07973_ (
  .A1(_02662_),
  .A2(\sresult[28][11] ),
  .ZN(_02699_)
);

NAND2_X1 _07974_ (
  .A1(_02651_),
  .A2(din_61[11]),
  .ZN(_02700_)
);

NAND2_X1 _07975_ (
  .A1(_02699_),
  .A2(_02700_),
  .ZN(_02701_)
);

NAND2_X1 _07976_ (
  .A1(_02701_),
  .A2(_02654_),
  .ZN(_02702_)
);

NAND2_X1 _07977_ (
  .A1(_02667_),
  .A2(\sresult[29][11] ),
  .ZN(_02703_)
);

NAND2_X1 _07978_ (
  .A1(_02702_),
  .A2(_02703_),
  .ZN(_00359_)
);

NAND2_X1 _07979_ (
  .A1(_02662_),
  .A2(\sresult[29][0] ),
  .ZN(_02704_)
);

BUF_X4 _07980_ (
  .A(_02650_),
  .Z(_02705_)
);

NAND2_X1 _07981_ (
  .A1(_02705_),
  .A2(din_52[0]),
  .ZN(_02706_)
);

NAND2_X1 _07982_ (
  .A1(_02704_),
  .A2(_02706_),
  .ZN(_02707_)
);

BUF_X2 _07983_ (
  .A(_02544_),
  .Z(_02708_)
);

NAND2_X1 _07984_ (
  .A1(_02707_),
  .A2(_02708_),
  .ZN(_02709_)
);

NAND2_X1 _07985_ (
  .A1(_02667_),
  .A2(\sresult[30][0] ),
  .ZN(_02710_)
);

NAND2_X1 _07986_ (
  .A1(_02709_),
  .A2(_02710_),
  .ZN(_00360_)
);

NAND2_X1 _07987_ (
  .A1(_02662_),
  .A2(\sresult[29][1] ),
  .ZN(_02711_)
);

NAND2_X1 _07988_ (
  .A1(_02705_),
  .A2(din_52[1]),
  .ZN(_02712_)
);

NAND2_X1 _07989_ (
  .A1(_02711_),
  .A2(_02712_),
  .ZN(_02713_)
);

NAND2_X1 _07990_ (
  .A1(_02713_),
  .A2(_02708_),
  .ZN(_02714_)
);

NAND2_X1 _07991_ (
  .A1(_02667_),
  .A2(\sresult[30][1] ),
  .ZN(_02715_)
);

NAND2_X1 _07992_ (
  .A1(_02714_),
  .A2(_02715_),
  .ZN(_00361_)
);

BUF_X4 _07993_ (
  .A(_00800_),
  .Z(_02716_)
);

NAND2_X1 _07994_ (
  .A1(_02716_),
  .A2(\sresult[29][2] ),
  .ZN(_02717_)
);

NAND2_X1 _07995_ (
  .A1(_02705_),
  .A2(din_52[2]),
  .ZN(_02718_)
);

NAND2_X1 _07996_ (
  .A1(_02717_),
  .A2(_02718_),
  .ZN(_02719_)
);

NAND2_X1 _07997_ (
  .A1(_02719_),
  .A2(_02708_),
  .ZN(_02720_)
);

BUF_X1 _07998_ (
  .A(_00811_),
  .Z(_02721_)
);

NAND2_X1 _07999_ (
  .A1(_02721_),
  .A2(\sresult[30][2] ),
  .ZN(_02722_)
);

NAND2_X1 _08000_ (
  .A1(_02720_),
  .A2(_02722_),
  .ZN(_00362_)
);

NAND2_X1 _08001_ (
  .A1(_02716_),
  .A2(\sresult[29][3] ),
  .ZN(_02723_)
);

NAND2_X1 _08002_ (
  .A1(_02705_),
  .A2(din_52[3]),
  .ZN(_02724_)
);

NAND2_X1 _08003_ (
  .A1(_02723_),
  .A2(_02724_),
  .ZN(_02725_)
);

NAND2_X1 _08004_ (
  .A1(_02725_),
  .A2(_02708_),
  .ZN(_02726_)
);

NAND2_X1 _08005_ (
  .A1(_02721_),
  .A2(\sresult[30][3] ),
  .ZN(_02727_)
);

NAND2_X1 _08006_ (
  .A1(_02726_),
  .A2(_02727_),
  .ZN(_00363_)
);

NAND2_X1 _08007_ (
  .A1(_02716_),
  .A2(\sresult[29][4] ),
  .ZN(_02728_)
);

NAND2_X1 _08008_ (
  .A1(_02705_),
  .A2(din_52[4]),
  .ZN(_02729_)
);

NAND2_X1 _08009_ (
  .A1(_02728_),
  .A2(_02729_),
  .ZN(_02730_)
);

NAND2_X1 _08010_ (
  .A1(_02730_),
  .A2(_02708_),
  .ZN(_02731_)
);

NAND2_X1 _08011_ (
  .A1(_02721_),
  .A2(\sresult[30][4] ),
  .ZN(_02732_)
);

NAND2_X1 _08012_ (
  .A1(_02731_),
  .A2(_02732_),
  .ZN(_00364_)
);

NAND2_X1 _08013_ (
  .A1(_02716_),
  .A2(\sresult[29][5] ),
  .ZN(_02733_)
);

NAND2_X1 _08014_ (
  .A1(_02705_),
  .A2(din_52[5]),
  .ZN(_02734_)
);

NAND2_X1 _08015_ (
  .A1(_02733_),
  .A2(_02734_),
  .ZN(_02735_)
);

NAND2_X1 _08016_ (
  .A1(_02735_),
  .A2(_02708_),
  .ZN(_02736_)
);

NAND2_X1 _08017_ (
  .A1(_02721_),
  .A2(\sresult[30][5] ),
  .ZN(_02737_)
);

NAND2_X1 _08018_ (
  .A1(_02736_),
  .A2(_02737_),
  .ZN(_00365_)
);

NAND2_X1 _08019_ (
  .A1(_02716_),
  .A2(\sresult[29][6] ),
  .ZN(_02738_)
);

NAND2_X1 _08020_ (
  .A1(_02705_),
  .A2(din_52[6]),
  .ZN(_02739_)
);

NAND2_X1 _08021_ (
  .A1(_02738_),
  .A2(_02739_),
  .ZN(_02740_)
);

NAND2_X1 _08022_ (
  .A1(_02740_),
  .A2(_02708_),
  .ZN(_02741_)
);

NAND2_X1 _08023_ (
  .A1(_02721_),
  .A2(\sresult[30][6] ),
  .ZN(_02742_)
);

NAND2_X1 _08024_ (
  .A1(_02741_),
  .A2(_02742_),
  .ZN(_00366_)
);

NAND2_X1 _08025_ (
  .A1(_02716_),
  .A2(\sresult[29][7] ),
  .ZN(_02743_)
);

NAND2_X1 _08026_ (
  .A1(_02705_),
  .A2(din_52[7]),
  .ZN(_02744_)
);

NAND2_X1 _08027_ (
  .A1(_02743_),
  .A2(_02744_),
  .ZN(_02745_)
);

NAND2_X1 _08028_ (
  .A1(_02745_),
  .A2(_02708_),
  .ZN(_02746_)
);

NAND2_X1 _08029_ (
  .A1(_02721_),
  .A2(\sresult[30][7] ),
  .ZN(_02747_)
);

NAND2_X1 _08030_ (
  .A1(_02746_),
  .A2(_02747_),
  .ZN(_00367_)
);

NAND2_X1 _08031_ (
  .A1(_02716_),
  .A2(\sresult[29][8] ),
  .ZN(_02748_)
);

NAND2_X1 _08032_ (
  .A1(_02705_),
  .A2(din_52[8]),
  .ZN(_02749_)
);

NAND2_X1 _08033_ (
  .A1(_02748_),
  .A2(_02749_),
  .ZN(_02750_)
);

NAND2_X1 _08034_ (
  .A1(_02750_),
  .A2(_02708_),
  .ZN(_02751_)
);

NAND2_X1 _08035_ (
  .A1(_02721_),
  .A2(\sresult[30][8] ),
  .ZN(_02752_)
);

NAND2_X1 _08036_ (
  .A1(_02751_),
  .A2(_02752_),
  .ZN(_00368_)
);

NAND2_X1 _08037_ (
  .A1(_02716_),
  .A2(\sresult[29][9] ),
  .ZN(_02753_)
);

NAND2_X1 _08038_ (
  .A1(_02705_),
  .A2(din_52[9]),
  .ZN(_02754_)
);

NAND2_X1 _08039_ (
  .A1(_02753_),
  .A2(_02754_),
  .ZN(_02755_)
);

NAND2_X1 _08040_ (
  .A1(_02755_),
  .A2(_02708_),
  .ZN(_02756_)
);

NAND2_X1 _08041_ (
  .A1(_02721_),
  .A2(\sresult[30][9] ),
  .ZN(_02757_)
);

NAND2_X1 _08042_ (
  .A1(_02756_),
  .A2(_02757_),
  .ZN(_00369_)
);

NAND2_X1 _08043_ (
  .A1(_02716_),
  .A2(\sresult[29][10] ),
  .ZN(_02758_)
);

BUF_X4 _08044_ (
  .A(_02650_),
  .Z(_02759_)
);

NAND2_X1 _08045_ (
  .A1(_02759_),
  .A2(din_52[10]),
  .ZN(_02760_)
);

NAND2_X1 _08046_ (
  .A1(_02758_),
  .A2(_02760_),
  .ZN(_02761_)
);

BUF_X2 _08047_ (
  .A(_02544_),
  .Z(_02762_)
);

NAND2_X1 _08048_ (
  .A1(_02761_),
  .A2(_02762_),
  .ZN(_02763_)
);

NAND2_X1 _08049_ (
  .A1(_02721_),
  .A2(\sresult[30][10] ),
  .ZN(_02764_)
);

NAND2_X1 _08050_ (
  .A1(_02763_),
  .A2(_02764_),
  .ZN(_00370_)
);

NAND2_X1 _08051_ (
  .A1(_02716_),
  .A2(\sresult[29][11] ),
  .ZN(_02765_)
);

NAND2_X1 _08052_ (
  .A1(_02759_),
  .A2(din_52[11]),
  .ZN(_02766_)
);

NAND2_X1 _08053_ (
  .A1(_02765_),
  .A2(_02766_),
  .ZN(_02767_)
);

NAND2_X1 _08054_ (
  .A1(_02767_),
  .A2(_02762_),
  .ZN(_02768_)
);

NAND2_X1 _08055_ (
  .A1(_02721_),
  .A2(\sresult[30][11] ),
  .ZN(_02769_)
);

NAND2_X1 _08056_ (
  .A1(_02768_),
  .A2(_02769_),
  .ZN(_00371_)
);

BUF_X4 _08057_ (
  .A(_00800_),
  .Z(_02770_)
);

NAND2_X1 _08058_ (
  .A1(_02770_),
  .A2(\sresult[30][0] ),
  .ZN(_02771_)
);

NAND2_X1 _08059_ (
  .A1(_02759_),
  .A2(din_43[0]),
  .ZN(_02772_)
);

NAND2_X1 _08060_ (
  .A1(_02771_),
  .A2(_02772_),
  .ZN(_02773_)
);

NAND2_X1 _08061_ (
  .A1(_02773_),
  .A2(_02762_),
  .ZN(_02774_)
);

BUF_X1 _08062_ (
  .A(_00811_),
  .Z(_02775_)
);

NAND2_X1 _08063_ (
  .A1(_02775_),
  .A2(\sresult[31][0] ),
  .ZN(_02776_)
);

NAND2_X1 _08064_ (
  .A1(_02774_),
  .A2(_02776_),
  .ZN(_00372_)
);

NAND2_X1 _08065_ (
  .A1(_02770_),
  .A2(\sresult[30][1] ),
  .ZN(_02777_)
);

NAND2_X1 _08066_ (
  .A1(_02759_),
  .A2(din_43[1]),
  .ZN(_02778_)
);

NAND2_X1 _08067_ (
  .A1(_02777_),
  .A2(_02778_),
  .ZN(_02779_)
);

NAND2_X1 _08068_ (
  .A1(_02779_),
  .A2(_02762_),
  .ZN(_02780_)
);

NAND2_X1 _08069_ (
  .A1(_02775_),
  .A2(\sresult[31][1] ),
  .ZN(_02781_)
);

NAND2_X1 _08070_ (
  .A1(_02780_),
  .A2(_02781_),
  .ZN(_00373_)
);

NAND2_X1 _08071_ (
  .A1(_02770_),
  .A2(\sresult[30][2] ),
  .ZN(_02782_)
);

NAND2_X1 _08072_ (
  .A1(_02759_),
  .A2(din_43[2]),
  .ZN(_02783_)
);

NAND2_X1 _08073_ (
  .A1(_02782_),
  .A2(_02783_),
  .ZN(_02784_)
);

NAND2_X1 _08074_ (
  .A1(_02784_),
  .A2(_02762_),
  .ZN(_02785_)
);

NAND2_X1 _08075_ (
  .A1(_02775_),
  .A2(\sresult[31][2] ),
  .ZN(_02786_)
);

NAND2_X1 _08076_ (
  .A1(_02785_),
  .A2(_02786_),
  .ZN(_00374_)
);

NAND2_X1 _08077_ (
  .A1(_02770_),
  .A2(\sresult[30][3] ),
  .ZN(_02787_)
);

NAND2_X1 _08078_ (
  .A1(_02759_),
  .A2(din_43[3]),
  .ZN(_02788_)
);

NAND2_X1 _08079_ (
  .A1(_02787_),
  .A2(_02788_),
  .ZN(_02789_)
);

NAND2_X1 _08080_ (
  .A1(_02789_),
  .A2(_02762_),
  .ZN(_02790_)
);

NAND2_X1 _08081_ (
  .A1(_02775_),
  .A2(\sresult[31][3] ),
  .ZN(_02791_)
);

NAND2_X1 _08082_ (
  .A1(_02790_),
  .A2(_02791_),
  .ZN(_00375_)
);

NAND2_X1 _08083_ (
  .A1(_02770_),
  .A2(\sresult[30][4] ),
  .ZN(_02792_)
);

NAND2_X1 _08084_ (
  .A1(_02759_),
  .A2(din_43[4]),
  .ZN(_02793_)
);

NAND2_X1 _08085_ (
  .A1(_02792_),
  .A2(_02793_),
  .ZN(_02794_)
);

NAND2_X1 _08086_ (
  .A1(_02794_),
  .A2(_02762_),
  .ZN(_02795_)
);

NAND2_X1 _08087_ (
  .A1(_02775_),
  .A2(\sresult[31][4] ),
  .ZN(_02796_)
);

NAND2_X1 _08088_ (
  .A1(_02795_),
  .A2(_02796_),
  .ZN(_00376_)
);

NAND2_X1 _08089_ (
  .A1(_02770_),
  .A2(\sresult[30][5] ),
  .ZN(_02797_)
);

NAND2_X1 _08090_ (
  .A1(_02759_),
  .A2(din_43[5]),
  .ZN(_02798_)
);

NAND2_X1 _08091_ (
  .A1(_02797_),
  .A2(_02798_),
  .ZN(_02799_)
);

NAND2_X1 _08092_ (
  .A1(_02799_),
  .A2(_02762_),
  .ZN(_02800_)
);

NAND2_X1 _08093_ (
  .A1(_02775_),
  .A2(\sresult[31][5] ),
  .ZN(_02801_)
);

NAND2_X1 _08094_ (
  .A1(_02800_),
  .A2(_02801_),
  .ZN(_00377_)
);

NAND2_X1 _08095_ (
  .A1(_02770_),
  .A2(\sresult[30][6] ),
  .ZN(_02802_)
);

NAND2_X1 _08096_ (
  .A1(_02759_),
  .A2(din_43[6]),
  .ZN(_02803_)
);

NAND2_X1 _08097_ (
  .A1(_02802_),
  .A2(_02803_),
  .ZN(_02804_)
);

NAND2_X1 _08098_ (
  .A1(_02804_),
  .A2(_02762_),
  .ZN(_02805_)
);

NAND2_X1 _08099_ (
  .A1(_02775_),
  .A2(\sresult[31][6] ),
  .ZN(_02806_)
);

NAND2_X1 _08100_ (
  .A1(_02805_),
  .A2(_02806_),
  .ZN(_00378_)
);

NAND2_X1 _08101_ (
  .A1(_02770_),
  .A2(\sresult[30][7] ),
  .ZN(_02807_)
);

NAND2_X1 _08102_ (
  .A1(_02759_),
  .A2(din_43[7]),
  .ZN(_02808_)
);

NAND2_X1 _08103_ (
  .A1(_02807_),
  .A2(_02808_),
  .ZN(_02809_)
);

NAND2_X1 _08104_ (
  .A1(_02809_),
  .A2(_02762_),
  .ZN(_02810_)
);

NAND2_X1 _08105_ (
  .A1(_02775_),
  .A2(\sresult[31][7] ),
  .ZN(_02811_)
);

NAND2_X1 _08106_ (
  .A1(_02810_),
  .A2(_02811_),
  .ZN(_00379_)
);

NAND2_X1 _08107_ (
  .A1(_02770_),
  .A2(\sresult[30][8] ),
  .ZN(_02812_)
);

BUF_X4 _08108_ (
  .A(_02650_),
  .Z(_02813_)
);

NAND2_X1 _08109_ (
  .A1(_02813_),
  .A2(din_43[8]),
  .ZN(_02814_)
);

NAND2_X1 _08110_ (
  .A1(_02812_),
  .A2(_02814_),
  .ZN(_02815_)
);

BUF_X2 _08111_ (
  .A(_02544_),
  .Z(_02816_)
);

NAND2_X1 _08112_ (
  .A1(_02815_),
  .A2(_02816_),
  .ZN(_02817_)
);

NAND2_X1 _08113_ (
  .A1(_02775_),
  .A2(\sresult[31][8] ),
  .ZN(_02818_)
);

NAND2_X1 _08114_ (
  .A1(_02817_),
  .A2(_02818_),
  .ZN(_00380_)
);

NAND2_X1 _08115_ (
  .A1(_02770_),
  .A2(\sresult[30][9] ),
  .ZN(_02819_)
);

NAND2_X1 _08116_ (
  .A1(_02813_),
  .A2(din_43[9]),
  .ZN(_02820_)
);

NAND2_X1 _08117_ (
  .A1(_02819_),
  .A2(_02820_),
  .ZN(_02821_)
);

NAND2_X1 _08118_ (
  .A1(_02821_),
  .A2(_02816_),
  .ZN(_02822_)
);

NAND2_X1 _08119_ (
  .A1(_02775_),
  .A2(\sresult[31][9] ),
  .ZN(_02823_)
);

NAND2_X1 _08120_ (
  .A1(_02822_),
  .A2(_02823_),
  .ZN(_00381_)
);

NAND2_X1 _08121_ (
  .A1(_00801_),
  .A2(\sresult[30][10] ),
  .ZN(_02824_)
);

NAND2_X1 _08122_ (
  .A1(_02813_),
  .A2(din_43[10]),
  .ZN(_02825_)
);

NAND2_X1 _08123_ (
  .A1(_02824_),
  .A2(_02825_),
  .ZN(_02826_)
);

NAND2_X1 _08124_ (
  .A1(_02826_),
  .A2(_02816_),
  .ZN(_02827_)
);

NAND2_X1 _08125_ (
  .A1(_00812_),
  .A2(\sresult[31][10] ),
  .ZN(_02828_)
);

NAND2_X1 _08126_ (
  .A1(_02827_),
  .A2(_02828_),
  .ZN(_00382_)
);

NAND2_X1 _08127_ (
  .A1(_00801_),
  .A2(\sresult[30][11] ),
  .ZN(_02829_)
);

NAND2_X1 _08128_ (
  .A1(_02813_),
  .A2(din_43[11]),
  .ZN(_02830_)
);

NAND2_X1 _08129_ (
  .A1(_02829_),
  .A2(_02830_),
  .ZN(_02831_)
);

NAND2_X1 _08130_ (
  .A1(_02831_),
  .A2(_02816_),
  .ZN(_02832_)
);

NAND2_X1 _08131_ (
  .A1(_00812_),
  .A2(\sresult[31][11] ),
  .ZN(_02833_)
);

NAND2_X1 _08132_ (
  .A1(_02832_),
  .A2(_02833_),
  .ZN(_00383_)
);

NAND2_X1 _08133_ (
  .A1(_00801_),
  .A2(\sresult[31][0] ),
  .ZN(_02834_)
);

NAND2_X1 _08134_ (
  .A1(_02813_),
  .A2(din_34[0]),
  .ZN(_02835_)
);

NAND2_X1 _08135_ (
  .A1(_02834_),
  .A2(_02835_),
  .ZN(_02836_)
);

NAND2_X1 _08136_ (
  .A1(_02836_),
  .A2(_02816_),
  .ZN(_02837_)
);

NAND2_X1 _08137_ (
  .A1(_00812_),
  .A2(\sresult[32][0] ),
  .ZN(_02838_)
);

NAND2_X1 _08138_ (
  .A1(_02837_),
  .A2(_02838_),
  .ZN(_00384_)
);

NAND2_X1 _08139_ (
  .A1(_00801_),
  .A2(\sresult[31][1] ),
  .ZN(_02839_)
);

NAND2_X1 _08140_ (
  .A1(_02813_),
  .A2(din_34[1]),
  .ZN(_02840_)
);

NAND2_X1 _08141_ (
  .A1(_02839_),
  .A2(_02840_),
  .ZN(_02841_)
);

NAND2_X1 _08142_ (
  .A1(_02841_),
  .A2(_02816_),
  .ZN(_02842_)
);

NAND2_X1 _08143_ (
  .A1(_00812_),
  .A2(\sresult[32][1] ),
  .ZN(_02843_)
);

NAND2_X1 _08144_ (
  .A1(_02842_),
  .A2(_02843_),
  .ZN(_00385_)
);

NAND2_X1 _08145_ (
  .A1(_00801_),
  .A2(\sresult[31][2] ),
  .ZN(_02844_)
);

NAND2_X1 _08146_ (
  .A1(_02813_),
  .A2(din_34[2]),
  .ZN(_02845_)
);

NAND2_X1 _08147_ (
  .A1(_02844_),
  .A2(_02845_),
  .ZN(_02846_)
);

NAND2_X1 _08148_ (
  .A1(_02846_),
  .A2(_02816_),
  .ZN(_02847_)
);

NAND2_X1 _08149_ (
  .A1(_00812_),
  .A2(\sresult[32][2] ),
  .ZN(_02848_)
);

NAND2_X1 _08150_ (
  .A1(_02847_),
  .A2(_02848_),
  .ZN(_00386_)
);

NAND2_X1 _08151_ (
  .A1(_00801_),
  .A2(\sresult[31][3] ),
  .ZN(_02849_)
);

NAND2_X1 _08152_ (
  .A1(_00803_),
  .A2(din_34[3]),
  .ZN(_02850_)
);

NAND2_X1 _08153_ (
  .A1(_02849_),
  .A2(_02850_),
  .ZN(_02851_)
);

NAND2_X1 _08154_ (
  .A1(_02851_),
  .A2(_02816_),
  .ZN(_02852_)
);

NAND2_X1 _08155_ (
  .A1(_00812_),
  .A2(\sresult[32][3] ),
  .ZN(_02853_)
);

NAND2_X1 _08156_ (
  .A1(_02852_),
  .A2(_02853_),
  .ZN(_00387_)
);

NAND2_X1 _08157_ (
  .A1(_00801_),
  .A2(\sresult[31][4] ),
  .ZN(_02854_)
);

NAND2_X1 _08158_ (
  .A1(_02813_),
  .A2(din_34[4]),
  .ZN(_02855_)
);

NAND2_X1 _08159_ (
  .A1(_02854_),
  .A2(_02855_),
  .ZN(_02856_)
);

NAND2_X1 _08160_ (
  .A1(_02856_),
  .A2(_00807_),
  .ZN(_02857_)
);

NAND2_X1 _08161_ (
  .A1(_00812_),
  .A2(\sresult[32][4] ),
  .ZN(_02858_)
);

NAND2_X1 _08162_ (
  .A1(_02857_),
  .A2(_02858_),
  .ZN(_00388_)
);

NAND2_X1 _08163_ (
  .A1(_00801_),
  .A2(\sresult[31][5] ),
  .ZN(_02859_)
);

NAND2_X1 _08164_ (
  .A1(_00803_),
  .A2(din_34[5]),
  .ZN(_02860_)
);

NAND2_X1 _08165_ (
  .A1(_02859_),
  .A2(_02860_),
  .ZN(_02861_)
);

NAND2_X1 _08166_ (
  .A1(_02861_),
  .A2(_02816_),
  .ZN(_02862_)
);

NAND2_X1 _08167_ (
  .A1(_00812_),
  .A2(\sresult[32][5] ),
  .ZN(_02863_)
);

NAND2_X1 _08168_ (
  .A1(_02862_),
  .A2(_02863_),
  .ZN(_00389_)
);

NAND2_X1 _08169_ (
  .A1(_00814_),
  .A2(\sresult[31][6] ),
  .ZN(_02864_)
);

BUF_X4 _08170_ (
  .A(_02650_),
  .Z(_02865_)
);

NAND2_X1 _08171_ (
  .A1(_02865_),
  .A2(din_34[6]),
  .ZN(_02866_)
);

NAND2_X1 _08172_ (
  .A1(_02864_),
  .A2(_02866_),
  .ZN(_02867_)
);

NAND2_X1 _08173_ (
  .A1(_02867_),
  .A2(_00807_),
  .ZN(_02868_)
);

NAND2_X1 _08174_ (
  .A1(_00820_),
  .A2(\sresult[32][6] ),
  .ZN(_02869_)
);

NAND2_X1 _08175_ (
  .A1(_02868_),
  .A2(_02869_),
  .ZN(_00390_)
);

NAND2_X1 _08176_ (
  .A1(_00801_),
  .A2(\sresult[31][7] ),
  .ZN(_02870_)
);

NAND2_X1 _08177_ (
  .A1(_02865_),
  .A2(din_34[7]),
  .ZN(_02871_)
);

NAND2_X1 _08178_ (
  .A1(_02870_),
  .A2(_02871_),
  .ZN(_02872_)
);

BUF_X2 _08179_ (
  .A(_02544_),
  .Z(_02873_)
);

NAND2_X1 _08180_ (
  .A1(_02872_),
  .A2(_02873_),
  .ZN(_02874_)
);

NAND2_X1 _08181_ (
  .A1(_00812_),
  .A2(\sresult[32][7] ),
  .ZN(_02875_)
);

NAND2_X1 _08182_ (
  .A1(_02874_),
  .A2(_02875_),
  .ZN(_00391_)
);

BUF_X4 _08183_ (
  .A(_00800_),
  .Z(_02876_)
);

NAND2_X1 _08184_ (
  .A1(_02876_),
  .A2(\sresult[31][8] ),
  .ZN(_02877_)
);

NAND2_X1 _08185_ (
  .A1(_02865_),
  .A2(din_34[8]),
  .ZN(_02878_)
);

NAND2_X1 _08186_ (
  .A1(_02877_),
  .A2(_02878_),
  .ZN(_02879_)
);

NAND2_X1 _08187_ (
  .A1(_02879_),
  .A2(_02873_),
  .ZN(_02880_)
);

BUF_X1 _08188_ (
  .A(_00811_),
  .Z(_02881_)
);

NAND2_X1 _08189_ (
  .A1(_02881_),
  .A2(\sresult[32][8] ),
  .ZN(_02882_)
);

NAND2_X1 _08190_ (
  .A1(_02880_),
  .A2(_02882_),
  .ZN(_00392_)
);

NAND2_X1 _08191_ (
  .A1(_02876_),
  .A2(\sresult[31][9] ),
  .ZN(_02883_)
);

NAND2_X1 _08192_ (
  .A1(_02865_),
  .A2(din_34[9]),
  .ZN(_02884_)
);

NAND2_X1 _08193_ (
  .A1(_02883_),
  .A2(_02884_),
  .ZN(_02885_)
);

NAND2_X1 _08194_ (
  .A1(_02885_),
  .A2(_02873_),
  .ZN(_02886_)
);

NAND2_X1 _08195_ (
  .A1(_02881_),
  .A2(\sresult[32][9] ),
  .ZN(_02887_)
);

NAND2_X1 _08196_ (
  .A1(_02886_),
  .A2(_02887_),
  .ZN(_00393_)
);

NAND2_X1 _08197_ (
  .A1(_02876_),
  .A2(\sresult[31][10] ),
  .ZN(_02888_)
);

NAND2_X1 _08198_ (
  .A1(_02865_),
  .A2(din_34[10]),
  .ZN(_02889_)
);

NAND2_X1 _08199_ (
  .A1(_02888_),
  .A2(_02889_),
  .ZN(_02890_)
);

NAND2_X1 _08200_ (
  .A1(_02890_),
  .A2(_02873_),
  .ZN(_02891_)
);

NAND2_X1 _08201_ (
  .A1(_02881_),
  .A2(\sresult[32][10] ),
  .ZN(_02892_)
);

NAND2_X1 _08202_ (
  .A1(_02891_),
  .A2(_02892_),
  .ZN(_00394_)
);

NAND2_X1 _08203_ (
  .A1(_02876_),
  .A2(\sresult[31][11] ),
  .ZN(_02893_)
);

NAND2_X1 _08204_ (
  .A1(_02865_),
  .A2(din_34[11]),
  .ZN(_02894_)
);

NAND2_X1 _08205_ (
  .A1(_02893_),
  .A2(_02894_),
  .ZN(_02895_)
);

NAND2_X1 _08206_ (
  .A1(_02895_),
  .A2(_02873_),
  .ZN(_02896_)
);

NAND2_X1 _08207_ (
  .A1(_02881_),
  .A2(\sresult[32][11] ),
  .ZN(_02897_)
);

NAND2_X1 _08208_ (
  .A1(_02896_),
  .A2(_02897_),
  .ZN(_00395_)
);

NAND2_X1 _08209_ (
  .A1(_02876_),
  .A2(\sresult[32][0] ),
  .ZN(_02898_)
);

NAND2_X1 _08210_ (
  .A1(_02865_),
  .A2(din_25[0]),
  .ZN(_02899_)
);

NAND2_X1 _08211_ (
  .A1(_02898_),
  .A2(_02899_),
  .ZN(_02900_)
);

NAND2_X1 _08212_ (
  .A1(_02900_),
  .A2(_02873_),
  .ZN(_02901_)
);

NAND2_X1 _08213_ (
  .A1(_02881_),
  .A2(\sresult[33][0] ),
  .ZN(_02902_)
);

NAND2_X1 _08214_ (
  .A1(_02901_),
  .A2(_02902_),
  .ZN(_00396_)
);

NAND2_X1 _08215_ (
  .A1(_02876_),
  .A2(\sresult[32][1] ),
  .ZN(_02903_)
);

NAND2_X1 _08216_ (
  .A1(_02865_),
  .A2(din_25[1]),
  .ZN(_02904_)
);

NAND2_X1 _08217_ (
  .A1(_02903_),
  .A2(_02904_),
  .ZN(_02905_)
);

NAND2_X1 _08218_ (
  .A1(_02905_),
  .A2(_02873_),
  .ZN(_02906_)
);

NAND2_X1 _08219_ (
  .A1(_02881_),
  .A2(\sresult[33][1] ),
  .ZN(_02907_)
);

NAND2_X1 _08220_ (
  .A1(_02906_),
  .A2(_02907_),
  .ZN(_00397_)
);

NAND2_X1 _08221_ (
  .A1(_02876_),
  .A2(\sresult[32][2] ),
  .ZN(_02908_)
);

NAND2_X1 _08222_ (
  .A1(_02865_),
  .A2(din_25[2]),
  .ZN(_02909_)
);

NAND2_X1 _08223_ (
  .A1(_02908_),
  .A2(_02909_),
  .ZN(_02910_)
);

NAND2_X1 _08224_ (
  .A1(_02910_),
  .A2(_02873_),
  .ZN(_02911_)
);

NAND2_X1 _08225_ (
  .A1(_02881_),
  .A2(\sresult[33][2] ),
  .ZN(_02912_)
);

NAND2_X1 _08226_ (
  .A1(_02911_),
  .A2(_02912_),
  .ZN(_00398_)
);

NAND2_X1 _08227_ (
  .A1(_02876_),
  .A2(\sresult[32][3] ),
  .ZN(_02913_)
);

NAND2_X1 _08228_ (
  .A1(_02865_),
  .A2(din_25[3]),
  .ZN(_02914_)
);

NAND2_X1 _08229_ (
  .A1(_02913_),
  .A2(_02914_),
  .ZN(_02915_)
);

NAND2_X1 _08230_ (
  .A1(_02915_),
  .A2(_02873_),
  .ZN(_02916_)
);

NAND2_X1 _08231_ (
  .A1(_02881_),
  .A2(\sresult[33][3] ),
  .ZN(_02917_)
);

NAND2_X1 _08232_ (
  .A1(_02916_),
  .A2(_02917_),
  .ZN(_00399_)
);

NAND2_X1 _08233_ (
  .A1(_02876_),
  .A2(\sresult[32][4] ),
  .ZN(_02918_)
);

BUF_X4 _08234_ (
  .A(_02650_),
  .Z(_02919_)
);

NAND2_X1 _08235_ (
  .A1(_02919_),
  .A2(din_25[4]),
  .ZN(_02920_)
);

NAND2_X1 _08236_ (
  .A1(_02918_),
  .A2(_02920_),
  .ZN(_02921_)
);

BUF_X2 _08237_ (
  .A(_02544_),
  .Z(_02922_)
);

NAND2_X1 _08238_ (
  .A1(_02921_),
  .A2(_02922_),
  .ZN(_02923_)
);

NAND2_X1 _08239_ (
  .A1(_02881_),
  .A2(\sresult[33][4] ),
  .ZN(_02924_)
);

NAND2_X1 _08240_ (
  .A1(_02923_),
  .A2(_02924_),
  .ZN(_00400_)
);

NAND2_X1 _08241_ (
  .A1(_02876_),
  .A2(\sresult[32][5] ),
  .ZN(_02925_)
);

NAND2_X1 _08242_ (
  .A1(_02919_),
  .A2(din_25[5]),
  .ZN(_02926_)
);

NAND2_X1 _08243_ (
  .A1(_02925_),
  .A2(_02926_),
  .ZN(_02927_)
);

NAND2_X1 _08244_ (
  .A1(_02927_),
  .A2(_02922_),
  .ZN(_02928_)
);

NAND2_X1 _08245_ (
  .A1(_02881_),
  .A2(\sresult[33][5] ),
  .ZN(_02929_)
);

NAND2_X1 _08246_ (
  .A1(_02928_),
  .A2(_02929_),
  .ZN(_00401_)
);

BUF_X4 _08247_ (
  .A(_00800_),
  .Z(_02930_)
);

NAND2_X1 _08248_ (
  .A1(_02930_),
  .A2(\sresult[32][6] ),
  .ZN(_02931_)
);

NAND2_X1 _08249_ (
  .A1(_02919_),
  .A2(din_25[6]),
  .ZN(_02932_)
);

NAND2_X1 _08250_ (
  .A1(_02931_),
  .A2(_02932_),
  .ZN(_02933_)
);

NAND2_X1 _08251_ (
  .A1(_02933_),
  .A2(_02922_),
  .ZN(_02934_)
);

BUF_X1 _08252_ (
  .A(_00811_),
  .Z(_02935_)
);

NAND2_X1 _08253_ (
  .A1(_02935_),
  .A2(\sresult[33][6] ),
  .ZN(_02936_)
);

NAND2_X1 _08254_ (
  .A1(_02934_),
  .A2(_02936_),
  .ZN(_00402_)
);

NAND2_X1 _08255_ (
  .A1(_02930_),
  .A2(\sresult[32][7] ),
  .ZN(_02937_)
);

NAND2_X1 _08256_ (
  .A1(_02919_),
  .A2(din_25[7]),
  .ZN(_02938_)
);

NAND2_X1 _08257_ (
  .A1(_02937_),
  .A2(_02938_),
  .ZN(_02939_)
);

NAND2_X1 _08258_ (
  .A1(_02939_),
  .A2(_02922_),
  .ZN(_02940_)
);

NAND2_X1 _08259_ (
  .A1(_02935_),
  .A2(\sresult[33][7] ),
  .ZN(_02941_)
);

NAND2_X1 _08260_ (
  .A1(_02940_),
  .A2(_02941_),
  .ZN(_00403_)
);

NAND2_X1 _08261_ (
  .A1(_02930_),
  .A2(\sresult[32][8] ),
  .ZN(_02942_)
);

NAND2_X1 _08262_ (
  .A1(_02919_),
  .A2(din_25[8]),
  .ZN(_02943_)
);

NAND2_X1 _08263_ (
  .A1(_02942_),
  .A2(_02943_),
  .ZN(_02944_)
);

NAND2_X1 _08264_ (
  .A1(_02944_),
  .A2(_02922_),
  .ZN(_02945_)
);

NAND2_X1 _08265_ (
  .A1(_02935_),
  .A2(\sresult[33][8] ),
  .ZN(_02946_)
);

NAND2_X1 _08266_ (
  .A1(_02945_),
  .A2(_02946_),
  .ZN(_00404_)
);

NAND2_X1 _08267_ (
  .A1(_02930_),
  .A2(\sresult[32][9] ),
  .ZN(_02947_)
);

NAND2_X1 _08268_ (
  .A1(_02919_),
  .A2(din_25[9]),
  .ZN(_02948_)
);

NAND2_X1 _08269_ (
  .A1(_02947_),
  .A2(_02948_),
  .ZN(_02949_)
);

NAND2_X1 _08270_ (
  .A1(_02949_),
  .A2(_02922_),
  .ZN(_02950_)
);

NAND2_X1 _08271_ (
  .A1(_02935_),
  .A2(\sresult[33][9] ),
  .ZN(_02951_)
);

NAND2_X1 _08272_ (
  .A1(_02950_),
  .A2(_02951_),
  .ZN(_00405_)
);

NAND2_X1 _08273_ (
  .A1(_02930_),
  .A2(\sresult[32][10] ),
  .ZN(_02952_)
);

NAND2_X1 _08274_ (
  .A1(_02919_),
  .A2(din_25[10]),
  .ZN(_02953_)
);

NAND2_X1 _08275_ (
  .A1(_02952_),
  .A2(_02953_),
  .ZN(_02954_)
);

NAND2_X1 _08276_ (
  .A1(_02954_),
  .A2(_02922_),
  .ZN(_02955_)
);

NAND2_X1 _08277_ (
  .A1(_02935_),
  .A2(\sresult[33][10] ),
  .ZN(_02956_)
);

NAND2_X1 _08278_ (
  .A1(_02955_),
  .A2(_02956_),
  .ZN(_00406_)
);

NAND2_X1 _08279_ (
  .A1(_02930_),
  .A2(\sresult[32][11] ),
  .ZN(_02957_)
);

NAND2_X1 _08280_ (
  .A1(_02919_),
  .A2(din_25[11]),
  .ZN(_02958_)
);

NAND2_X1 _08281_ (
  .A1(_02957_),
  .A2(_02958_),
  .ZN(_02959_)
);

NAND2_X1 _08282_ (
  .A1(_02959_),
  .A2(_02922_),
  .ZN(_02960_)
);

NAND2_X1 _08283_ (
  .A1(_02935_),
  .A2(\sresult[33][11] ),
  .ZN(_02961_)
);

NAND2_X1 _08284_ (
  .A1(_02960_),
  .A2(_02961_),
  .ZN(_00407_)
);

NAND2_X1 _08285_ (
  .A1(_02930_),
  .A2(\sresult[33][0] ),
  .ZN(_02962_)
);

NAND2_X1 _08286_ (
  .A1(_02919_),
  .A2(din_16[0]),
  .ZN(_02963_)
);

NAND2_X1 _08287_ (
  .A1(_02962_),
  .A2(_02963_),
  .ZN(_02964_)
);

NAND2_X1 _08288_ (
  .A1(_02964_),
  .A2(_02922_),
  .ZN(_02965_)
);

NAND2_X1 _08289_ (
  .A1(_02935_),
  .A2(\sresult[34][0] ),
  .ZN(_02966_)
);

NAND2_X1 _08290_ (
  .A1(_02965_),
  .A2(_02966_),
  .ZN(_00408_)
);

NAND2_X1 _08291_ (
  .A1(_02930_),
  .A2(\sresult[33][1] ),
  .ZN(_02967_)
);

NAND2_X1 _08292_ (
  .A1(_02919_),
  .A2(din_16[1]),
  .ZN(_02968_)
);

NAND2_X1 _08293_ (
  .A1(_02967_),
  .A2(_02968_),
  .ZN(_02969_)
);

NAND2_X1 _08294_ (
  .A1(_02969_),
  .A2(_02922_),
  .ZN(_02970_)
);

NAND2_X1 _08295_ (
  .A1(_02935_),
  .A2(\sresult[34][1] ),
  .ZN(_02971_)
);

NAND2_X1 _08296_ (
  .A1(_02970_),
  .A2(_02971_),
  .ZN(_00409_)
);

NAND2_X1 _08297_ (
  .A1(_02930_),
  .A2(\sresult[33][2] ),
  .ZN(_02972_)
);

BUF_X4 _08298_ (
  .A(_02650_),
  .Z(_02973_)
);

NAND2_X1 _08299_ (
  .A1(_02973_),
  .A2(din_16[2]),
  .ZN(_02974_)
);

NAND2_X1 _08300_ (
  .A1(_02972_),
  .A2(_02974_),
  .ZN(_02975_)
);

BUF_X2 _08301_ (
  .A(_02544_),
  .Z(_02976_)
);

NAND2_X1 _08302_ (
  .A1(_02975_),
  .A2(_02976_),
  .ZN(_02977_)
);

NAND2_X1 _08303_ (
  .A1(_02935_),
  .A2(\sresult[34][2] ),
  .ZN(_02978_)
);

NAND2_X1 _08304_ (
  .A1(_02977_),
  .A2(_02978_),
  .ZN(_00410_)
);

NAND2_X1 _08305_ (
  .A1(_02930_),
  .A2(\sresult[33][3] ),
  .ZN(_02979_)
);

NAND2_X1 _08306_ (
  .A1(_02973_),
  .A2(din_16[3]),
  .ZN(_02980_)
);

NAND2_X1 _08307_ (
  .A1(_02979_),
  .A2(_02980_),
  .ZN(_02981_)
);

NAND2_X1 _08308_ (
  .A1(_02981_),
  .A2(_02976_),
  .ZN(_02982_)
);

NAND2_X1 _08309_ (
  .A1(_02935_),
  .A2(\sresult[34][3] ),
  .ZN(_02983_)
);

NAND2_X1 _08310_ (
  .A1(_02982_),
  .A2(_02983_),
  .ZN(_00411_)
);

BUF_X4 _08311_ (
  .A(_00800_),
  .Z(_02984_)
);

NAND2_X1 _08312_ (
  .A1(_02984_),
  .A2(\sresult[33][4] ),
  .ZN(_02985_)
);

NAND2_X1 _08313_ (
  .A1(_02973_),
  .A2(din_16[4]),
  .ZN(_02986_)
);

NAND2_X1 _08314_ (
  .A1(_02985_),
  .A2(_02986_),
  .ZN(_02987_)
);

NAND2_X1 _08315_ (
  .A1(_02987_),
  .A2(_02976_),
  .ZN(_02988_)
);

BUF_X1 _08316_ (
  .A(_00811_),
  .Z(_02989_)
);

NAND2_X1 _08317_ (
  .A1(_02989_),
  .A2(\sresult[34][4] ),
  .ZN(_02990_)
);

NAND2_X1 _08318_ (
  .A1(_02988_),
  .A2(_02990_),
  .ZN(_00412_)
);

NAND2_X1 _08319_ (
  .A1(_02984_),
  .A2(\sresult[33][5] ),
  .ZN(_02991_)
);

NAND2_X1 _08320_ (
  .A1(_02973_),
  .A2(din_16[5]),
  .ZN(_02992_)
);

NAND2_X1 _08321_ (
  .A1(_02991_),
  .A2(_02992_),
  .ZN(_02993_)
);

NAND2_X1 _08322_ (
  .A1(_02993_),
  .A2(_02976_),
  .ZN(_02994_)
);

NAND2_X1 _08323_ (
  .A1(_02989_),
  .A2(\sresult[34][5] ),
  .ZN(_02995_)
);

NAND2_X1 _08324_ (
  .A1(_02994_),
  .A2(_02995_),
  .ZN(_00413_)
);

NAND2_X1 _08325_ (
  .A1(_02984_),
  .A2(\sresult[33][6] ),
  .ZN(_02996_)
);

NAND2_X1 _08326_ (
  .A1(_02973_),
  .A2(din_16[6]),
  .ZN(_02997_)
);

NAND2_X1 _08327_ (
  .A1(_02996_),
  .A2(_02997_),
  .ZN(_02998_)
);

NAND2_X1 _08328_ (
  .A1(_02998_),
  .A2(_02976_),
  .ZN(_02999_)
);

NAND2_X1 _08329_ (
  .A1(_02989_),
  .A2(\sresult[34][6] ),
  .ZN(_03000_)
);

NAND2_X1 _08330_ (
  .A1(_02999_),
  .A2(_03000_),
  .ZN(_00414_)
);

NAND2_X1 _08331_ (
  .A1(_02984_),
  .A2(\sresult[33][7] ),
  .ZN(_03001_)
);

NAND2_X1 _08332_ (
  .A1(_02973_),
  .A2(din_16[7]),
  .ZN(_03002_)
);

NAND2_X1 _08333_ (
  .A1(_03001_),
  .A2(_03002_),
  .ZN(_03003_)
);

NAND2_X1 _08334_ (
  .A1(_03003_),
  .A2(_02976_),
  .ZN(_03004_)
);

NAND2_X1 _08335_ (
  .A1(_02989_),
  .A2(\sresult[34][7] ),
  .ZN(_03005_)
);

NAND2_X1 _08336_ (
  .A1(_03004_),
  .A2(_03005_),
  .ZN(_00415_)
);

NAND2_X1 _08337_ (
  .A1(_02984_),
  .A2(\sresult[33][8] ),
  .ZN(_03006_)
);

NAND2_X1 _08338_ (
  .A1(_02973_),
  .A2(din_16[8]),
  .ZN(_03007_)
);

NAND2_X1 _08339_ (
  .A1(_03006_),
  .A2(_03007_),
  .ZN(_03008_)
);

NAND2_X1 _08340_ (
  .A1(_03008_),
  .A2(_02976_),
  .ZN(_03009_)
);

NAND2_X1 _08341_ (
  .A1(_02989_),
  .A2(\sresult[34][8] ),
  .ZN(_03010_)
);

NAND2_X1 _08342_ (
  .A1(_03009_),
  .A2(_03010_),
  .ZN(_00416_)
);

NAND2_X1 _08343_ (
  .A1(_02984_),
  .A2(\sresult[33][9] ),
  .ZN(_03011_)
);

NAND2_X1 _08344_ (
  .A1(_02973_),
  .A2(din_16[9]),
  .ZN(_03012_)
);

NAND2_X1 _08345_ (
  .A1(_03011_),
  .A2(_03012_),
  .ZN(_03013_)
);

NAND2_X1 _08346_ (
  .A1(_03013_),
  .A2(_02976_),
  .ZN(_03014_)
);

NAND2_X1 _08347_ (
  .A1(_02989_),
  .A2(\sresult[34][9] ),
  .ZN(_03015_)
);

NAND2_X1 _08348_ (
  .A1(_03014_),
  .A2(_03015_),
  .ZN(_00417_)
);

NAND2_X1 _08349_ (
  .A1(_02984_),
  .A2(\sresult[33][10] ),
  .ZN(_03016_)
);

NAND2_X1 _08350_ (
  .A1(_02973_),
  .A2(din_16[10]),
  .ZN(_03017_)
);

NAND2_X1 _08351_ (
  .A1(_03016_),
  .A2(_03017_),
  .ZN(_03018_)
);

NAND2_X1 _08352_ (
  .A1(_03018_),
  .A2(_02976_),
  .ZN(_03019_)
);

NAND2_X1 _08353_ (
  .A1(_02989_),
  .A2(\sresult[34][10] ),
  .ZN(_03020_)
);

NAND2_X1 _08354_ (
  .A1(_03019_),
  .A2(_03020_),
  .ZN(_00418_)
);

NAND2_X1 _08355_ (
  .A1(_02984_),
  .A2(\sresult[33][11] ),
  .ZN(_03021_)
);

NAND2_X1 _08356_ (
  .A1(_02973_),
  .A2(din_16[11]),
  .ZN(_03022_)
);

NAND2_X1 _08357_ (
  .A1(_03021_),
  .A2(_03022_),
  .ZN(_03023_)
);

NAND2_X1 _08358_ (
  .A1(_03023_),
  .A2(_02976_),
  .ZN(_03024_)
);

NAND2_X1 _08359_ (
  .A1(_02989_),
  .A2(\sresult[34][11] ),
  .ZN(_03025_)
);

NAND2_X1 _08360_ (
  .A1(_03024_),
  .A2(_03025_),
  .ZN(_00419_)
);

NAND2_X1 _08361_ (
  .A1(_02984_),
  .A2(\sresult[34][0] ),
  .ZN(_03026_)
);

BUF_X4 _08362_ (
  .A(_02650_),
  .Z(_03027_)
);

NAND2_X1 _08363_ (
  .A1(_03027_),
  .A2(din_07[0]),
  .ZN(_03028_)
);

NAND2_X1 _08364_ (
  .A1(_03026_),
  .A2(_03028_),
  .ZN(_03029_)
);

BUF_X2 _08365_ (
  .A(_02544_),
  .Z(_03030_)
);

NAND2_X1 _08366_ (
  .A1(_03029_),
  .A2(_03030_),
  .ZN(_03031_)
);

NAND2_X1 _08367_ (
  .A1(_02989_),
  .A2(\sresult[35][0] ),
  .ZN(_03032_)
);

NAND2_X1 _08368_ (
  .A1(_03031_),
  .A2(_03032_),
  .ZN(_00420_)
);

NAND2_X1 _08369_ (
  .A1(_02984_),
  .A2(\sresult[34][1] ),
  .ZN(_03033_)
);

NAND2_X1 _08370_ (
  .A1(_03027_),
  .A2(din_07[1]),
  .ZN(_03034_)
);

NAND2_X1 _08371_ (
  .A1(_03033_),
  .A2(_03034_),
  .ZN(_03035_)
);

NAND2_X1 _08372_ (
  .A1(_03035_),
  .A2(_03030_),
  .ZN(_03036_)
);

NAND2_X1 _08373_ (
  .A1(_02989_),
  .A2(\sresult[35][1] ),
  .ZN(_03037_)
);

NAND2_X1 _08374_ (
  .A1(_03036_),
  .A2(_03037_),
  .ZN(_00421_)
);

BUF_X4 _08375_ (
  .A(_00800_),
  .Z(_03038_)
);

NAND2_X1 _08376_ (
  .A1(_03038_),
  .A2(\sresult[34][2] ),
  .ZN(_03039_)
);

NAND2_X1 _08377_ (
  .A1(_03027_),
  .A2(din_07[2]),
  .ZN(_03040_)
);

NAND2_X1 _08378_ (
  .A1(_03039_),
  .A2(_03040_),
  .ZN(_03041_)
);

NAND2_X1 _08379_ (
  .A1(_03041_),
  .A2(_03030_),
  .ZN(_03042_)
);

BUF_X1 _08380_ (
  .A(_00811_),
  .Z(_03043_)
);

NAND2_X1 _08381_ (
  .A1(_03043_),
  .A2(\sresult[35][2] ),
  .ZN(_03044_)
);

NAND2_X1 _08382_ (
  .A1(_03042_),
  .A2(_03044_),
  .ZN(_00422_)
);

NAND2_X1 _08383_ (
  .A1(_03038_),
  .A2(\sresult[34][3] ),
  .ZN(_03045_)
);

NAND2_X1 _08384_ (
  .A1(_03027_),
  .A2(din_07[3]),
  .ZN(_03046_)
);

NAND2_X1 _08385_ (
  .A1(_03045_),
  .A2(_03046_),
  .ZN(_03047_)
);

NAND2_X1 _08386_ (
  .A1(_03047_),
  .A2(_03030_),
  .ZN(_03048_)
);

NAND2_X1 _08387_ (
  .A1(_03043_),
  .A2(\sresult[35][3] ),
  .ZN(_03049_)
);

NAND2_X1 _08388_ (
  .A1(_03048_),
  .A2(_03049_),
  .ZN(_00423_)
);

NAND2_X1 _08389_ (
  .A1(_03038_),
  .A2(\sresult[34][4] ),
  .ZN(_03050_)
);

NAND2_X1 _08390_ (
  .A1(_03027_),
  .A2(din_07[4]),
  .ZN(_03051_)
);

NAND2_X1 _08391_ (
  .A1(_03050_),
  .A2(_03051_),
  .ZN(_03052_)
);

NAND2_X1 _08392_ (
  .A1(_03052_),
  .A2(_03030_),
  .ZN(_03053_)
);

NAND2_X1 _08393_ (
  .A1(_03043_),
  .A2(\sresult[35][4] ),
  .ZN(_03054_)
);

NAND2_X1 _08394_ (
  .A1(_03053_),
  .A2(_03054_),
  .ZN(_00424_)
);

NAND2_X1 _08395_ (
  .A1(_03038_),
  .A2(\sresult[34][5] ),
  .ZN(_03055_)
);

NAND2_X1 _08396_ (
  .A1(_03027_),
  .A2(din_07[5]),
  .ZN(_03056_)
);

NAND2_X1 _08397_ (
  .A1(_03055_),
  .A2(_03056_),
  .ZN(_03057_)
);

NAND2_X1 _08398_ (
  .A1(_03057_),
  .A2(_03030_),
  .ZN(_03058_)
);

NAND2_X1 _08399_ (
  .A1(_03043_),
  .A2(\sresult[35][5] ),
  .ZN(_03059_)
);

NAND2_X1 _08400_ (
  .A1(_03058_),
  .A2(_03059_),
  .ZN(_00425_)
);

NAND2_X1 _08401_ (
  .A1(_03038_),
  .A2(\sresult[34][6] ),
  .ZN(_03060_)
);

NAND2_X1 _08402_ (
  .A1(_03027_),
  .A2(din_07[6]),
  .ZN(_03061_)
);

NAND2_X1 _08403_ (
  .A1(_03060_),
  .A2(_03061_),
  .ZN(_03062_)
);

NAND2_X1 _08404_ (
  .A1(_03062_),
  .A2(_03030_),
  .ZN(_03063_)
);

NAND2_X1 _08405_ (
  .A1(_03043_),
  .A2(\sresult[35][6] ),
  .ZN(_03064_)
);

NAND2_X1 _08406_ (
  .A1(_03063_),
  .A2(_03064_),
  .ZN(_00426_)
);

NAND2_X1 _08407_ (
  .A1(_03038_),
  .A2(\sresult[34][7] ),
  .ZN(_03065_)
);

NAND2_X1 _08408_ (
  .A1(_03027_),
  .A2(din_07[7]),
  .ZN(_03066_)
);

NAND2_X1 _08409_ (
  .A1(_03065_),
  .A2(_03066_),
  .ZN(_03067_)
);

NAND2_X1 _08410_ (
  .A1(_03067_),
  .A2(_03030_),
  .ZN(_03068_)
);

NAND2_X1 _08411_ (
  .A1(_03043_),
  .A2(\sresult[35][7] ),
  .ZN(_03069_)
);

NAND2_X1 _08412_ (
  .A1(_03068_),
  .A2(_03069_),
  .ZN(_00427_)
);

NAND2_X1 _08413_ (
  .A1(_03038_),
  .A2(\sresult[34][8] ),
  .ZN(_03070_)
);

NAND2_X1 _08414_ (
  .A1(_03027_),
  .A2(din_07[8]),
  .ZN(_03071_)
);

NAND2_X1 _08415_ (
  .A1(_03070_),
  .A2(_03071_),
  .ZN(_03072_)
);

NAND2_X1 _08416_ (
  .A1(_03072_),
  .A2(_03030_),
  .ZN(_03073_)
);

NAND2_X1 _08417_ (
  .A1(_03043_),
  .A2(\sresult[35][8] ),
  .ZN(_03074_)
);

NAND2_X1 _08418_ (
  .A1(_03073_),
  .A2(_03074_),
  .ZN(_00428_)
);

NAND2_X1 _08419_ (
  .A1(_03038_),
  .A2(\sresult[34][9] ),
  .ZN(_03075_)
);

NAND2_X1 _08420_ (
  .A1(_03027_),
  .A2(din_07[9]),
  .ZN(_03076_)
);

NAND2_X1 _08421_ (
  .A1(_03075_),
  .A2(_03076_),
  .ZN(_03077_)
);

NAND2_X1 _08422_ (
  .A1(_03077_),
  .A2(_03030_),
  .ZN(_03078_)
);

NAND2_X1 _08423_ (
  .A1(_03043_),
  .A2(\sresult[35][9] ),
  .ZN(_03079_)
);

NAND2_X1 _08424_ (
  .A1(_03078_),
  .A2(_03079_),
  .ZN(_00429_)
);

NAND2_X1 _08425_ (
  .A1(_03038_),
  .A2(\sresult[34][10] ),
  .ZN(_03080_)
);

BUF_X4 _08426_ (
  .A(_02650_),
  .Z(_03081_)
);

NAND2_X1 _08427_ (
  .A1(_03081_),
  .A2(din_07[10]),
  .ZN(_03082_)
);

NAND2_X1 _08428_ (
  .A1(_03080_),
  .A2(_03082_),
  .ZN(_03083_)
);

BUF_X4 _08429_ (
  .A(_00911_),
  .Z(_03084_)
);

BUF_X2 _08430_ (
  .A(_03084_),
  .Z(_03085_)
);

NAND2_X1 _08431_ (
  .A1(_03083_),
  .A2(_03085_),
  .ZN(_03086_)
);

NAND2_X1 _08432_ (
  .A1(_03043_),
  .A2(\sresult[35][10] ),
  .ZN(_03087_)
);

NAND2_X1 _08433_ (
  .A1(_03086_),
  .A2(_03087_),
  .ZN(_00430_)
);

NAND2_X1 _08434_ (
  .A1(_03038_),
  .A2(\sresult[34][11] ),
  .ZN(_03088_)
);

NAND2_X1 _08435_ (
  .A1(_03081_),
  .A2(din_07[11]),
  .ZN(_03089_)
);

NAND2_X1 _08436_ (
  .A1(_03088_),
  .A2(_03089_),
  .ZN(_03090_)
);

NAND2_X1 _08437_ (
  .A1(_03090_),
  .A2(_03085_),
  .ZN(_03091_)
);

NAND2_X1 _08438_ (
  .A1(_03043_),
  .A2(\sresult[35][11] ),
  .ZN(_03092_)
);

NAND2_X1 _08439_ (
  .A1(_03091_),
  .A2(_03092_),
  .ZN(_00431_)
);

BUF_X4 _08440_ (
  .A(_00800_),
  .Z(_03093_)
);

NAND2_X1 _08441_ (
  .A1(_03093_),
  .A2(\sresult[35][0] ),
  .ZN(_03094_)
);

NAND2_X1 _08442_ (
  .A1(_03081_),
  .A2(din_06[0]),
  .ZN(_03095_)
);

NAND2_X1 _08443_ (
  .A1(_03094_),
  .A2(_03095_),
  .ZN(_03096_)
);

NAND2_X1 _08444_ (
  .A1(_03096_),
  .A2(_03085_),
  .ZN(_03097_)
);

BUF_X1 _08445_ (
  .A(_00811_),
  .Z(_03098_)
);

NAND2_X1 _08446_ (
  .A1(_03098_),
  .A2(\sresult[36][0] ),
  .ZN(_03099_)
);

NAND2_X1 _08447_ (
  .A1(_03097_),
  .A2(_03099_),
  .ZN(_00432_)
);

NAND2_X1 _08448_ (
  .A1(_03093_),
  .A2(\sresult[35][1] ),
  .ZN(_03100_)
);

NAND2_X1 _08449_ (
  .A1(_03081_),
  .A2(din_06[1]),
  .ZN(_03101_)
);

NAND2_X1 _08450_ (
  .A1(_03100_),
  .A2(_03101_),
  .ZN(_03102_)
);

NAND2_X1 _08451_ (
  .A1(_03102_),
  .A2(_03085_),
  .ZN(_03103_)
);

NAND2_X1 _08452_ (
  .A1(_03098_),
  .A2(\sresult[36][1] ),
  .ZN(_03104_)
);

NAND2_X1 _08453_ (
  .A1(_03103_),
  .A2(_03104_),
  .ZN(_00433_)
);

NAND2_X1 _08454_ (
  .A1(_03093_),
  .A2(\sresult[35][2] ),
  .ZN(_03105_)
);

NAND2_X1 _08455_ (
  .A1(_03081_),
  .A2(din_06[2]),
  .ZN(_03106_)
);

NAND2_X1 _08456_ (
  .A1(_03105_),
  .A2(_03106_),
  .ZN(_03107_)
);

NAND2_X1 _08457_ (
  .A1(_03107_),
  .A2(_03085_),
  .ZN(_03108_)
);

NAND2_X1 _08458_ (
  .A1(_03098_),
  .A2(\sresult[36][2] ),
  .ZN(_03109_)
);

NAND2_X1 _08459_ (
  .A1(_03108_),
  .A2(_03109_),
  .ZN(_00434_)
);

NAND2_X1 _08460_ (
  .A1(_03093_),
  .A2(\sresult[35][3] ),
  .ZN(_03110_)
);

NAND2_X1 _08461_ (
  .A1(_03081_),
  .A2(din_06[3]),
  .ZN(_03111_)
);

NAND2_X1 _08462_ (
  .A1(_03110_),
  .A2(_03111_),
  .ZN(_03112_)
);

NAND2_X1 _08463_ (
  .A1(_03112_),
  .A2(_03085_),
  .ZN(_03113_)
);

NAND2_X1 _08464_ (
  .A1(_03098_),
  .A2(\sresult[36][3] ),
  .ZN(_03114_)
);

NAND2_X1 _08465_ (
  .A1(_03113_),
  .A2(_03114_),
  .ZN(_00435_)
);

NAND2_X1 _08466_ (
  .A1(_03093_),
  .A2(\sresult[35][4] ),
  .ZN(_03115_)
);

NAND2_X1 _08467_ (
  .A1(_03081_),
  .A2(din_06[4]),
  .ZN(_03116_)
);

NAND2_X1 _08468_ (
  .A1(_03115_),
  .A2(_03116_),
  .ZN(_03117_)
);

NAND2_X1 _08469_ (
  .A1(_03117_),
  .A2(_03085_),
  .ZN(_03118_)
);

NAND2_X1 _08470_ (
  .A1(_03098_),
  .A2(\sresult[36][4] ),
  .ZN(_03119_)
);

NAND2_X1 _08471_ (
  .A1(_03118_),
  .A2(_03119_),
  .ZN(_00436_)
);

NAND2_X1 _08472_ (
  .A1(_03093_),
  .A2(\sresult[35][5] ),
  .ZN(_03120_)
);

NAND2_X1 _08473_ (
  .A1(_03081_),
  .A2(din_06[5]),
  .ZN(_03121_)
);

NAND2_X1 _08474_ (
  .A1(_03120_),
  .A2(_03121_),
  .ZN(_03122_)
);

NAND2_X1 _08475_ (
  .A1(_03122_),
  .A2(_03085_),
  .ZN(_03123_)
);

NAND2_X1 _08476_ (
  .A1(_03098_),
  .A2(\sresult[36][5] ),
  .ZN(_03124_)
);

NAND2_X1 _08477_ (
  .A1(_03123_),
  .A2(_03124_),
  .ZN(_00437_)
);

NAND2_X1 _08478_ (
  .A1(_03093_),
  .A2(\sresult[35][6] ),
  .ZN(_03125_)
);

NAND2_X1 _08479_ (
  .A1(_03081_),
  .A2(din_06[6]),
  .ZN(_03126_)
);

NAND2_X1 _08480_ (
  .A1(_03125_),
  .A2(_03126_),
  .ZN(_03127_)
);

NAND2_X1 _08481_ (
  .A1(_03127_),
  .A2(_03085_),
  .ZN(_03128_)
);

NAND2_X1 _08482_ (
  .A1(_03098_),
  .A2(\sresult[36][6] ),
  .ZN(_03129_)
);

NAND2_X1 _08483_ (
  .A1(_03128_),
  .A2(_03129_),
  .ZN(_00438_)
);

NAND2_X1 _08484_ (
  .A1(_03093_),
  .A2(\sresult[35][7] ),
  .ZN(_03130_)
);

NAND2_X1 _08485_ (
  .A1(_03081_),
  .A2(din_06[7]),
  .ZN(_03131_)
);

NAND2_X1 _08486_ (
  .A1(_03130_),
  .A2(_03131_),
  .ZN(_03132_)
);

NAND2_X1 _08487_ (
  .A1(_03132_),
  .A2(_03085_),
  .ZN(_03133_)
);

NAND2_X1 _08488_ (
  .A1(_03098_),
  .A2(\sresult[36][7] ),
  .ZN(_03134_)
);

NAND2_X1 _08489_ (
  .A1(_03133_),
  .A2(_03134_),
  .ZN(_00439_)
);

NAND2_X1 _08490_ (
  .A1(_03093_),
  .A2(\sresult[35][8] ),
  .ZN(_03135_)
);

BUF_X4 _08491_ (
  .A(_02650_),
  .Z(_03136_)
);

NAND2_X1 _08492_ (
  .A1(_03136_),
  .A2(din_06[8]),
  .ZN(_03137_)
);

NAND2_X1 _08493_ (
  .A1(_03135_),
  .A2(_03137_),
  .ZN(_03138_)
);

BUF_X2 _08494_ (
  .A(_03084_),
  .Z(_03139_)
);

NAND2_X1 _08495_ (
  .A1(_03138_),
  .A2(_03139_),
  .ZN(_03140_)
);

NAND2_X1 _08496_ (
  .A1(_03098_),
  .A2(\sresult[36][8] ),
  .ZN(_03141_)
);

NAND2_X1 _08497_ (
  .A1(_03140_),
  .A2(_03141_),
  .ZN(_00440_)
);

NAND2_X1 _08498_ (
  .A1(_03093_),
  .A2(\sresult[35][9] ),
  .ZN(_03142_)
);

NAND2_X1 _08499_ (
  .A1(_03136_),
  .A2(din_06[9]),
  .ZN(_03143_)
);

NAND2_X1 _08500_ (
  .A1(_03142_),
  .A2(_03143_),
  .ZN(_03144_)
);

NAND2_X1 _08501_ (
  .A1(_03144_),
  .A2(_03139_),
  .ZN(_03145_)
);

NAND2_X1 _08502_ (
  .A1(_03098_),
  .A2(\sresult[36][9] ),
  .ZN(_03146_)
);

NAND2_X1 _08503_ (
  .A1(_03145_),
  .A2(_03146_),
  .ZN(_00441_)
);

BUF_X8 _08504_ (
  .A(_00799_),
  .Z(_03147_)
);

BUF_X4 _08505_ (
  .A(_03147_),
  .Z(_03148_)
);

NAND2_X1 _08506_ (
  .A1(_03148_),
  .A2(\sresult[35][10] ),
  .ZN(_03149_)
);

NAND2_X1 _08507_ (
  .A1(_03136_),
  .A2(din_06[10]),
  .ZN(_03150_)
);

NAND2_X1 _08508_ (
  .A1(_03149_),
  .A2(_03150_),
  .ZN(_03151_)
);

NAND2_X1 _08509_ (
  .A1(_03151_),
  .A2(_03139_),
  .ZN(_03152_)
);

BUF_X1 _08510_ (
  .A(_00811_),
  .Z(_03153_)
);

NAND2_X1 _08511_ (
  .A1(_03153_),
  .A2(\sresult[36][10] ),
  .ZN(_03154_)
);

NAND2_X1 _08512_ (
  .A1(_03152_),
  .A2(_03154_),
  .ZN(_00442_)
);

NAND2_X1 _08513_ (
  .A1(_03148_),
  .A2(\sresult[35][11] ),
  .ZN(_03155_)
);

NAND2_X1 _08514_ (
  .A1(_03136_),
  .A2(din_06[11]),
  .ZN(_03156_)
);

NAND2_X1 _08515_ (
  .A1(_03155_),
  .A2(_03156_),
  .ZN(_03157_)
);

NAND2_X1 _08516_ (
  .A1(_03157_),
  .A2(_03139_),
  .ZN(_03158_)
);

NAND2_X1 _08517_ (
  .A1(_03153_),
  .A2(\sresult[36][11] ),
  .ZN(_03159_)
);

NAND2_X1 _08518_ (
  .A1(_03158_),
  .A2(_03159_),
  .ZN(_00443_)
);

NAND2_X1 _08519_ (
  .A1(_03148_),
  .A2(\sresult[36][0] ),
  .ZN(_03160_)
);

NAND2_X1 _08520_ (
  .A1(_03136_),
  .A2(din_15[0]),
  .ZN(_03161_)
);

NAND2_X1 _08521_ (
  .A1(_03160_),
  .A2(_03161_),
  .ZN(_03162_)
);

NAND2_X1 _08522_ (
  .A1(_03162_),
  .A2(_03139_),
  .ZN(_03163_)
);

NAND2_X1 _08523_ (
  .A1(_03153_),
  .A2(\sresult[37][0] ),
  .ZN(_03164_)
);

NAND2_X1 _08524_ (
  .A1(_03163_),
  .A2(_03164_),
  .ZN(_00444_)
);

NAND2_X1 _08525_ (
  .A1(_03148_),
  .A2(\sresult[36][1] ),
  .ZN(_03165_)
);

NAND2_X1 _08526_ (
  .A1(_03136_),
  .A2(din_15[1]),
  .ZN(_03166_)
);

NAND2_X1 _08527_ (
  .A1(_03165_),
  .A2(_03166_),
  .ZN(_03167_)
);

NAND2_X1 _08528_ (
  .A1(_03167_),
  .A2(_03139_),
  .ZN(_03168_)
);

NAND2_X1 _08529_ (
  .A1(_03153_),
  .A2(\sresult[37][1] ),
  .ZN(_03169_)
);

NAND2_X1 _08530_ (
  .A1(_03168_),
  .A2(_03169_),
  .ZN(_00445_)
);

NAND2_X1 _08531_ (
  .A1(_03148_),
  .A2(\sresult[36][2] ),
  .ZN(_03170_)
);

NAND2_X1 _08532_ (
  .A1(_03136_),
  .A2(din_15[2]),
  .ZN(_03171_)
);

NAND2_X1 _08533_ (
  .A1(_03170_),
  .A2(_03171_),
  .ZN(_03172_)
);

NAND2_X1 _08534_ (
  .A1(_03172_),
  .A2(_03139_),
  .ZN(_03173_)
);

NAND2_X1 _08535_ (
  .A1(_03153_),
  .A2(\sresult[37][2] ),
  .ZN(_03174_)
);

NAND2_X1 _08536_ (
  .A1(_03173_),
  .A2(_03174_),
  .ZN(_00446_)
);

NAND2_X1 _08537_ (
  .A1(_03148_),
  .A2(\sresult[36][3] ),
  .ZN(_03175_)
);

NAND2_X1 _08538_ (
  .A1(_03136_),
  .A2(din_15[3]),
  .ZN(_03176_)
);

NAND2_X1 _08539_ (
  .A1(_03175_),
  .A2(_03176_),
  .ZN(_03177_)
);

NAND2_X1 _08540_ (
  .A1(_03177_),
  .A2(_03139_),
  .ZN(_03178_)
);

NAND2_X1 _08541_ (
  .A1(_03153_),
  .A2(\sresult[37][3] ),
  .ZN(_03179_)
);

NAND2_X1 _08542_ (
  .A1(_03178_),
  .A2(_03179_),
  .ZN(_00447_)
);

NAND2_X1 _08543_ (
  .A1(_03148_),
  .A2(\sresult[36][4] ),
  .ZN(_03180_)
);

NAND2_X1 _08544_ (
  .A1(_03136_),
  .A2(din_15[4]),
  .ZN(_03181_)
);

NAND2_X1 _08545_ (
  .A1(_03180_),
  .A2(_03181_),
  .ZN(_03182_)
);

NAND2_X1 _08546_ (
  .A1(_03182_),
  .A2(_03139_),
  .ZN(_03183_)
);

NAND2_X1 _08547_ (
  .A1(_03153_),
  .A2(\sresult[37][4] ),
  .ZN(_03184_)
);

NAND2_X1 _08548_ (
  .A1(_03183_),
  .A2(_03184_),
  .ZN(_00448_)
);

NAND2_X1 _08549_ (
  .A1(_03148_),
  .A2(\sresult[36][5] ),
  .ZN(_03185_)
);

NAND2_X1 _08550_ (
  .A1(_03136_),
  .A2(din_15[5]),
  .ZN(_03186_)
);

NAND2_X1 _08551_ (
  .A1(_03185_),
  .A2(_03186_),
  .ZN(_03187_)
);

NAND2_X1 _08552_ (
  .A1(_03187_),
  .A2(_03139_),
  .ZN(_03188_)
);

NAND2_X1 _08553_ (
  .A1(_03153_),
  .A2(\sresult[37][5] ),
  .ZN(_03189_)
);

NAND2_X1 _08554_ (
  .A1(_03188_),
  .A2(_03189_),
  .ZN(_00449_)
);

NAND2_X1 _08555_ (
  .A1(_03148_),
  .A2(\sresult[36][6] ),
  .ZN(_03190_)
);

BUF_X8 _08556_ (
  .A(_00770_),
  .Z(_03191_)
);

BUF_X4 _08557_ (
  .A(_03191_),
  .Z(_03192_)
);

NAND2_X1 _08558_ (
  .A1(_03192_),
  .A2(din_15[6]),
  .ZN(_03193_)
);

NAND2_X1 _08559_ (
  .A1(_03190_),
  .A2(_03193_),
  .ZN(_03194_)
);

BUF_X2 _08560_ (
  .A(_03084_),
  .Z(_03195_)
);

NAND2_X1 _08561_ (
  .A1(_03194_),
  .A2(_03195_),
  .ZN(_03196_)
);

NAND2_X1 _08562_ (
  .A1(_03153_),
  .A2(\sresult[37][6] ),
  .ZN(_03197_)
);

NAND2_X1 _08563_ (
  .A1(_03196_),
  .A2(_03197_),
  .ZN(_00450_)
);

NAND2_X1 _08564_ (
  .A1(_03148_),
  .A2(\sresult[36][7] ),
  .ZN(_03198_)
);

NAND2_X1 _08565_ (
  .A1(_03192_),
  .A2(din_15[7]),
  .ZN(_03199_)
);

NAND2_X1 _08566_ (
  .A1(_03198_),
  .A2(_03199_),
  .ZN(_03200_)
);

NAND2_X1 _08567_ (
  .A1(_03200_),
  .A2(_03195_),
  .ZN(_03201_)
);

NAND2_X1 _08568_ (
  .A1(_03153_),
  .A2(\sresult[37][7] ),
  .ZN(_03202_)
);

NAND2_X1 _08569_ (
  .A1(_03201_),
  .A2(_03202_),
  .ZN(_00451_)
);

BUF_X4 _08570_ (
  .A(_03147_),
  .Z(_03203_)
);

NAND2_X1 _08571_ (
  .A1(_03203_),
  .A2(\sresult[36][8] ),
  .ZN(_03204_)
);

NAND2_X1 _08572_ (
  .A1(_03192_),
  .A2(din_15[8]),
  .ZN(_03205_)
);

NAND2_X1 _08573_ (
  .A1(_03204_),
  .A2(_03205_),
  .ZN(_03206_)
);

NAND2_X1 _08574_ (
  .A1(_03206_),
  .A2(_03195_),
  .ZN(_03207_)
);

BUF_X8 _08575_ (
  .A(_00810_),
  .Z(_03208_)
);

BUF_X1 _08576_ (
  .A(_03208_),
  .Z(_03209_)
);

NAND2_X1 _08577_ (
  .A1(_03209_),
  .A2(\sresult[37][8] ),
  .ZN(_03210_)
);

NAND2_X1 _08578_ (
  .A1(_03207_),
  .A2(_03210_),
  .ZN(_00452_)
);

NAND2_X1 _08579_ (
  .A1(_03203_),
  .A2(\sresult[36][9] ),
  .ZN(_03211_)
);

NAND2_X1 _08580_ (
  .A1(_03192_),
  .A2(din_15[9]),
  .ZN(_03212_)
);

NAND2_X1 _08581_ (
  .A1(_03211_),
  .A2(_03212_),
  .ZN(_03213_)
);

NAND2_X1 _08582_ (
  .A1(_03213_),
  .A2(_03195_),
  .ZN(_03214_)
);

NAND2_X1 _08583_ (
  .A1(_03209_),
  .A2(\sresult[37][9] ),
  .ZN(_03215_)
);

NAND2_X1 _08584_ (
  .A1(_03214_),
  .A2(_03215_),
  .ZN(_00453_)
);

NAND2_X1 _08585_ (
  .A1(_03203_),
  .A2(\sresult[36][10] ),
  .ZN(_03216_)
);

NAND2_X1 _08586_ (
  .A1(_03192_),
  .A2(din_15[10]),
  .ZN(_03217_)
);

NAND2_X1 _08587_ (
  .A1(_03216_),
  .A2(_03217_),
  .ZN(_03218_)
);

NAND2_X1 _08588_ (
  .A1(_03218_),
  .A2(_03195_),
  .ZN(_03219_)
);

NAND2_X1 _08589_ (
  .A1(_03209_),
  .A2(\sresult[37][10] ),
  .ZN(_03220_)
);

NAND2_X1 _08590_ (
  .A1(_03219_),
  .A2(_03220_),
  .ZN(_00454_)
);

NAND2_X1 _08591_ (
  .A1(_03203_),
  .A2(\sresult[36][11] ),
  .ZN(_03221_)
);

NAND2_X1 _08592_ (
  .A1(_03192_),
  .A2(din_15[11]),
  .ZN(_03222_)
);

NAND2_X1 _08593_ (
  .A1(_03221_),
  .A2(_03222_),
  .ZN(_03223_)
);

NAND2_X1 _08594_ (
  .A1(_03223_),
  .A2(_03195_),
  .ZN(_03224_)
);

NAND2_X1 _08595_ (
  .A1(_03209_),
  .A2(\sresult[37][11] ),
  .ZN(_03225_)
);

NAND2_X1 _08596_ (
  .A1(_03224_),
  .A2(_03225_),
  .ZN(_00455_)
);

NAND2_X1 _08597_ (
  .A1(_03203_),
  .A2(\sresult[37][0] ),
  .ZN(_03226_)
);

NAND2_X1 _08598_ (
  .A1(_03192_),
  .A2(din_24[0]),
  .ZN(_03227_)
);

NAND2_X1 _08599_ (
  .A1(_03226_),
  .A2(_03227_),
  .ZN(_03228_)
);

NAND2_X1 _08600_ (
  .A1(_03228_),
  .A2(_03195_),
  .ZN(_03229_)
);

NAND2_X1 _08601_ (
  .A1(_03209_),
  .A2(\sresult[38][0] ),
  .ZN(_03230_)
);

NAND2_X1 _08602_ (
  .A1(_03229_),
  .A2(_03230_),
  .ZN(_00456_)
);

NAND2_X1 _08603_ (
  .A1(_03203_),
  .A2(\sresult[37][1] ),
  .ZN(_03231_)
);

NAND2_X1 _08604_ (
  .A1(_03192_),
  .A2(din_24[1]),
  .ZN(_03232_)
);

NAND2_X1 _08605_ (
  .A1(_03231_),
  .A2(_03232_),
  .ZN(_03233_)
);

NAND2_X1 _08606_ (
  .A1(_03233_),
  .A2(_03195_),
  .ZN(_03234_)
);

NAND2_X1 _08607_ (
  .A1(_03209_),
  .A2(\sresult[38][1] ),
  .ZN(_03235_)
);

NAND2_X1 _08608_ (
  .A1(_03234_),
  .A2(_03235_),
  .ZN(_00457_)
);

NAND2_X1 _08609_ (
  .A1(_03203_),
  .A2(\sresult[37][2] ),
  .ZN(_03236_)
);

NAND2_X1 _08610_ (
  .A1(_03192_),
  .A2(din_24[2]),
  .ZN(_03237_)
);

NAND2_X1 _08611_ (
  .A1(_03236_),
  .A2(_03237_),
  .ZN(_03238_)
);

NAND2_X1 _08612_ (
  .A1(_03238_),
  .A2(_03195_),
  .ZN(_03239_)
);

NAND2_X1 _08613_ (
  .A1(_03209_),
  .A2(\sresult[38][2] ),
  .ZN(_03240_)
);

NAND2_X1 _08614_ (
  .A1(_03239_),
  .A2(_03240_),
  .ZN(_00458_)
);

NAND2_X1 _08615_ (
  .A1(_03203_),
  .A2(\sresult[37][3] ),
  .ZN(_03241_)
);

NAND2_X1 _08616_ (
  .A1(_03192_),
  .A2(din_24[3]),
  .ZN(_03242_)
);

NAND2_X1 _08617_ (
  .A1(_03241_),
  .A2(_03242_),
  .ZN(_03243_)
);

NAND2_X1 _08618_ (
  .A1(_03243_),
  .A2(_03195_),
  .ZN(_03244_)
);

NAND2_X1 _08619_ (
  .A1(_03209_),
  .A2(\sresult[38][3] ),
  .ZN(_03245_)
);

NAND2_X1 _08620_ (
  .A1(_03244_),
  .A2(_03245_),
  .ZN(_00459_)
);

NAND2_X1 _08621_ (
  .A1(_03203_),
  .A2(\sresult[37][4] ),
  .ZN(_03246_)
);

BUF_X4 _08622_ (
  .A(_03191_),
  .Z(_03247_)
);

NAND2_X1 _08623_ (
  .A1(_03247_),
  .A2(din_24[4]),
  .ZN(_03248_)
);

NAND2_X1 _08624_ (
  .A1(_03246_),
  .A2(_03248_),
  .ZN(_03249_)
);

BUF_X2 _08625_ (
  .A(_03084_),
  .Z(_03250_)
);

NAND2_X1 _08626_ (
  .A1(_03249_),
  .A2(_03250_),
  .ZN(_03251_)
);

NAND2_X1 _08627_ (
  .A1(_03209_),
  .A2(\sresult[38][4] ),
  .ZN(_03252_)
);

NAND2_X1 _08628_ (
  .A1(_03251_),
  .A2(_03252_),
  .ZN(_00460_)
);

NAND2_X1 _08629_ (
  .A1(_03203_),
  .A2(\sresult[37][5] ),
  .ZN(_03253_)
);

NAND2_X1 _08630_ (
  .A1(_03247_),
  .A2(din_24[5]),
  .ZN(_03254_)
);

NAND2_X1 _08631_ (
  .A1(_03253_),
  .A2(_03254_),
  .ZN(_03255_)
);

NAND2_X1 _08632_ (
  .A1(_03255_),
  .A2(_03250_),
  .ZN(_03256_)
);

NAND2_X1 _08633_ (
  .A1(_03209_),
  .A2(\sresult[38][5] ),
  .ZN(_03257_)
);

NAND2_X1 _08634_ (
  .A1(_03256_),
  .A2(_03257_),
  .ZN(_00461_)
);

BUF_X4 _08635_ (
  .A(_03147_),
  .Z(_03258_)
);

NAND2_X1 _08636_ (
  .A1(_03258_),
  .A2(\sresult[37][6] ),
  .ZN(_03259_)
);

NAND2_X1 _08637_ (
  .A1(_03247_),
  .A2(din_24[6]),
  .ZN(_03260_)
);

NAND2_X1 _08638_ (
  .A1(_03259_),
  .A2(_03260_),
  .ZN(_03261_)
);

NAND2_X1 _08639_ (
  .A1(_03261_),
  .A2(_03250_),
  .ZN(_03262_)
);

BUF_X1 _08640_ (
  .A(_03208_),
  .Z(_03263_)
);

NAND2_X1 _08641_ (
  .A1(_03263_),
  .A2(\sresult[38][6] ),
  .ZN(_03264_)
);

NAND2_X1 _08642_ (
  .A1(_03262_),
  .A2(_03264_),
  .ZN(_00462_)
);

NAND2_X1 _08643_ (
  .A1(_03258_),
  .A2(\sresult[37][7] ),
  .ZN(_03265_)
);

NAND2_X1 _08644_ (
  .A1(_03247_),
  .A2(din_24[7]),
  .ZN(_03266_)
);

NAND2_X1 _08645_ (
  .A1(_03265_),
  .A2(_03266_),
  .ZN(_03267_)
);

NAND2_X1 _08646_ (
  .A1(_03267_),
  .A2(_03250_),
  .ZN(_03268_)
);

NAND2_X1 _08647_ (
  .A1(_03263_),
  .A2(\sresult[38][7] ),
  .ZN(_03269_)
);

NAND2_X1 _08648_ (
  .A1(_03268_),
  .A2(_03269_),
  .ZN(_00463_)
);

NAND2_X1 _08649_ (
  .A1(_03258_),
  .A2(\sresult[37][8] ),
  .ZN(_03270_)
);

NAND2_X1 _08650_ (
  .A1(_03247_),
  .A2(din_24[8]),
  .ZN(_03271_)
);

NAND2_X1 _08651_ (
  .A1(_03270_),
  .A2(_03271_),
  .ZN(_03272_)
);

NAND2_X1 _08652_ (
  .A1(_03272_),
  .A2(_03250_),
  .ZN(_03273_)
);

NAND2_X1 _08653_ (
  .A1(_03263_),
  .A2(\sresult[38][8] ),
  .ZN(_03274_)
);

NAND2_X1 _08654_ (
  .A1(_03273_),
  .A2(_03274_),
  .ZN(_00464_)
);

NAND2_X1 _08655_ (
  .A1(_03258_),
  .A2(\sresult[37][9] ),
  .ZN(_03275_)
);

NAND2_X1 _08656_ (
  .A1(_03247_),
  .A2(din_24[9]),
  .ZN(_03276_)
);

NAND2_X1 _08657_ (
  .A1(_03275_),
  .A2(_03276_),
  .ZN(_03277_)
);

NAND2_X1 _08658_ (
  .A1(_03277_),
  .A2(_03250_),
  .ZN(_03278_)
);

NAND2_X1 _08659_ (
  .A1(_03263_),
  .A2(\sresult[38][9] ),
  .ZN(_03279_)
);

NAND2_X1 _08660_ (
  .A1(_03278_),
  .A2(_03279_),
  .ZN(_00465_)
);

NAND2_X1 _08661_ (
  .A1(_03258_),
  .A2(\sresult[37][10] ),
  .ZN(_03280_)
);

NAND2_X1 _08662_ (
  .A1(_03247_),
  .A2(din_24[10]),
  .ZN(_03281_)
);

NAND2_X1 _08663_ (
  .A1(_03280_),
  .A2(_03281_),
  .ZN(_03282_)
);

NAND2_X1 _08664_ (
  .A1(_03282_),
  .A2(_03250_),
  .ZN(_03283_)
);

NAND2_X1 _08665_ (
  .A1(_03263_),
  .A2(\sresult[38][10] ),
  .ZN(_03284_)
);

NAND2_X1 _08666_ (
  .A1(_03283_),
  .A2(_03284_),
  .ZN(_00466_)
);

NAND2_X1 _08667_ (
  .A1(_03258_),
  .A2(\sresult[37][11] ),
  .ZN(_03285_)
);

NAND2_X1 _08668_ (
  .A1(_03247_),
  .A2(din_24[11]),
  .ZN(_03286_)
);

NAND2_X1 _08669_ (
  .A1(_03285_),
  .A2(_03286_),
  .ZN(_03287_)
);

NAND2_X1 _08670_ (
  .A1(_03287_),
  .A2(_03250_),
  .ZN(_03288_)
);

NAND2_X1 _08671_ (
  .A1(_03263_),
  .A2(\sresult[38][11] ),
  .ZN(_03289_)
);

NAND2_X1 _08672_ (
  .A1(_03288_),
  .A2(_03289_),
  .ZN(_00467_)
);

NAND2_X1 _08673_ (
  .A1(_03258_),
  .A2(\sresult[38][0] ),
  .ZN(_03290_)
);

NAND2_X1 _08674_ (
  .A1(_03247_),
  .A2(din_33[0]),
  .ZN(_03291_)
);

NAND2_X1 _08675_ (
  .A1(_03290_),
  .A2(_03291_),
  .ZN(_03292_)
);

NAND2_X1 _08676_ (
  .A1(_03292_),
  .A2(_03250_),
  .ZN(_03293_)
);

NAND2_X1 _08677_ (
  .A1(_03263_),
  .A2(\sresult[39][0] ),
  .ZN(_03294_)
);

NAND2_X1 _08678_ (
  .A1(_03293_),
  .A2(_03294_),
  .ZN(_00468_)
);

NAND2_X1 _08679_ (
  .A1(_03258_),
  .A2(\sresult[38][1] ),
  .ZN(_03295_)
);

NAND2_X1 _08680_ (
  .A1(_03247_),
  .A2(din_33[1]),
  .ZN(_03296_)
);

NAND2_X1 _08681_ (
  .A1(_03295_),
  .A2(_03296_),
  .ZN(_03297_)
);

NAND2_X1 _08682_ (
  .A1(_03297_),
  .A2(_03250_),
  .ZN(_03298_)
);

NAND2_X1 _08683_ (
  .A1(_03263_),
  .A2(\sresult[39][1] ),
  .ZN(_03299_)
);

NAND2_X1 _08684_ (
  .A1(_03298_),
  .A2(_03299_),
  .ZN(_00469_)
);

NAND2_X1 _08685_ (
  .A1(_03258_),
  .A2(\sresult[38][2] ),
  .ZN(_03300_)
);

BUF_X4 _08686_ (
  .A(_03191_),
  .Z(_03301_)
);

NAND2_X1 _08687_ (
  .A1(_03301_),
  .A2(din_33[2]),
  .ZN(_03302_)
);

NAND2_X1 _08688_ (
  .A1(_03300_),
  .A2(_03302_),
  .ZN(_03303_)
);

BUF_X2 _08689_ (
  .A(_03084_),
  .Z(_03304_)
);

NAND2_X1 _08690_ (
  .A1(_03303_),
  .A2(_03304_),
  .ZN(_03305_)
);

NAND2_X1 _08691_ (
  .A1(_03263_),
  .A2(\sresult[39][2] ),
  .ZN(_03306_)
);

NAND2_X1 _08692_ (
  .A1(_03305_),
  .A2(_03306_),
  .ZN(_00470_)
);

NAND2_X1 _08693_ (
  .A1(_03258_),
  .A2(\sresult[38][3] ),
  .ZN(_03307_)
);

NAND2_X1 _08694_ (
  .A1(_03301_),
  .A2(din_33[3]),
  .ZN(_03308_)
);

NAND2_X1 _08695_ (
  .A1(_03307_),
  .A2(_03308_),
  .ZN(_03309_)
);

NAND2_X1 _08696_ (
  .A1(_03309_),
  .A2(_03304_),
  .ZN(_03310_)
);

NAND2_X1 _08697_ (
  .A1(_03263_),
  .A2(\sresult[39][3] ),
  .ZN(_03311_)
);

NAND2_X1 _08698_ (
  .A1(_03310_),
  .A2(_03311_),
  .ZN(_00471_)
);

BUF_X4 _08699_ (
  .A(_03147_),
  .Z(_03312_)
);

NAND2_X1 _08700_ (
  .A1(_03312_),
  .A2(\sresult[38][4] ),
  .ZN(_03313_)
);

NAND2_X1 _08701_ (
  .A1(_03301_),
  .A2(din_33[4]),
  .ZN(_03314_)
);

NAND2_X1 _08702_ (
  .A1(_03313_),
  .A2(_03314_),
  .ZN(_03315_)
);

NAND2_X1 _08703_ (
  .A1(_03315_),
  .A2(_03304_),
  .ZN(_03316_)
);

BUF_X1 _08704_ (
  .A(_03208_),
  .Z(_03317_)
);

NAND2_X1 _08705_ (
  .A1(_03317_),
  .A2(\sresult[39][4] ),
  .ZN(_03318_)
);

NAND2_X1 _08706_ (
  .A1(_03316_),
  .A2(_03318_),
  .ZN(_00472_)
);

NAND2_X1 _08707_ (
  .A1(_03312_),
  .A2(\sresult[38][5] ),
  .ZN(_03319_)
);

NAND2_X1 _08708_ (
  .A1(_03301_),
  .A2(din_33[5]),
  .ZN(_03320_)
);

NAND2_X1 _08709_ (
  .A1(_03319_),
  .A2(_03320_),
  .ZN(_03321_)
);

NAND2_X1 _08710_ (
  .A1(_03321_),
  .A2(_03304_),
  .ZN(_03322_)
);

NAND2_X1 _08711_ (
  .A1(_03317_),
  .A2(\sresult[39][5] ),
  .ZN(_03323_)
);

NAND2_X1 _08712_ (
  .A1(_03322_),
  .A2(_03323_),
  .ZN(_00473_)
);

NAND2_X1 _08713_ (
  .A1(_03312_),
  .A2(\sresult[38][6] ),
  .ZN(_03324_)
);

NAND2_X1 _08714_ (
  .A1(_03301_),
  .A2(din_33[6]),
  .ZN(_03325_)
);

NAND2_X1 _08715_ (
  .A1(_03324_),
  .A2(_03325_),
  .ZN(_03326_)
);

NAND2_X1 _08716_ (
  .A1(_03326_),
  .A2(_03304_),
  .ZN(_03327_)
);

NAND2_X1 _08717_ (
  .A1(_03317_),
  .A2(\sresult[39][6] ),
  .ZN(_03328_)
);

NAND2_X1 _08718_ (
  .A1(_03327_),
  .A2(_03328_),
  .ZN(_00474_)
);

NAND2_X1 _08719_ (
  .A1(_03312_),
  .A2(\sresult[38][7] ),
  .ZN(_03329_)
);

NAND2_X1 _08720_ (
  .A1(_03301_),
  .A2(din_33[7]),
  .ZN(_03330_)
);

NAND2_X1 _08721_ (
  .A1(_03329_),
  .A2(_03330_),
  .ZN(_03331_)
);

NAND2_X1 _08722_ (
  .A1(_03331_),
  .A2(_03304_),
  .ZN(_03332_)
);

NAND2_X1 _08723_ (
  .A1(_03317_),
  .A2(\sresult[39][7] ),
  .ZN(_03333_)
);

NAND2_X1 _08724_ (
  .A1(_03332_),
  .A2(_03333_),
  .ZN(_00475_)
);

NAND2_X1 _08725_ (
  .A1(_03312_),
  .A2(\sresult[38][8] ),
  .ZN(_03334_)
);

NAND2_X1 _08726_ (
  .A1(_03301_),
  .A2(din_33[8]),
  .ZN(_03335_)
);

NAND2_X1 _08727_ (
  .A1(_03334_),
  .A2(_03335_),
  .ZN(_03336_)
);

NAND2_X1 _08728_ (
  .A1(_03336_),
  .A2(_03304_),
  .ZN(_03337_)
);

NAND2_X1 _08729_ (
  .A1(_03317_),
  .A2(\sresult[39][8] ),
  .ZN(_03338_)
);

NAND2_X1 _08730_ (
  .A1(_03337_),
  .A2(_03338_),
  .ZN(_00476_)
);

NAND2_X1 _08731_ (
  .A1(_03312_),
  .A2(\sresult[38][9] ),
  .ZN(_03339_)
);

NAND2_X1 _08732_ (
  .A1(_03301_),
  .A2(din_33[9]),
  .ZN(_03340_)
);

NAND2_X1 _08733_ (
  .A1(_03339_),
  .A2(_03340_),
  .ZN(_03341_)
);

NAND2_X1 _08734_ (
  .A1(_03341_),
  .A2(_03304_),
  .ZN(_03342_)
);

NAND2_X1 _08735_ (
  .A1(_03317_),
  .A2(\sresult[39][9] ),
  .ZN(_03343_)
);

NAND2_X1 _08736_ (
  .A1(_03342_),
  .A2(_03343_),
  .ZN(_00477_)
);

NAND2_X1 _08737_ (
  .A1(_03312_),
  .A2(\sresult[38][10] ),
  .ZN(_03344_)
);

NAND2_X1 _08738_ (
  .A1(_03301_),
  .A2(din_33[10]),
  .ZN(_03345_)
);

NAND2_X1 _08739_ (
  .A1(_03344_),
  .A2(_03345_),
  .ZN(_03346_)
);

NAND2_X1 _08740_ (
  .A1(_03346_),
  .A2(_03304_),
  .ZN(_03347_)
);

NAND2_X1 _08741_ (
  .A1(_03317_),
  .A2(\sresult[39][10] ),
  .ZN(_03348_)
);

NAND2_X1 _08742_ (
  .A1(_03347_),
  .A2(_03348_),
  .ZN(_00478_)
);

NAND2_X1 _08743_ (
  .A1(_03312_),
  .A2(\sresult[38][11] ),
  .ZN(_03349_)
);

NAND2_X1 _08744_ (
  .A1(_03301_),
  .A2(din_33[11]),
  .ZN(_03350_)
);

NAND2_X1 _08745_ (
  .A1(_03349_),
  .A2(_03350_),
  .ZN(_03351_)
);

NAND2_X1 _08746_ (
  .A1(_03351_),
  .A2(_03304_),
  .ZN(_03352_)
);

NAND2_X1 _08747_ (
  .A1(_03317_),
  .A2(\sresult[39][11] ),
  .ZN(_03353_)
);

NAND2_X1 _08748_ (
  .A1(_03352_),
  .A2(_03353_),
  .ZN(_00479_)
);

NAND2_X1 _08749_ (
  .A1(_03312_),
  .A2(\sresult[39][0] ),
  .ZN(_03354_)
);

BUF_X4 _08750_ (
  .A(_03191_),
  .Z(_03355_)
);

NAND2_X1 _08751_ (
  .A1(_03355_),
  .A2(din_42[0]),
  .ZN(_03356_)
);

NAND2_X1 _08752_ (
  .A1(_03354_),
  .A2(_03356_),
  .ZN(_03357_)
);

BUF_X2 _08753_ (
  .A(_03084_),
  .Z(_03358_)
);

NAND2_X1 _08754_ (
  .A1(_03357_),
  .A2(_03358_),
  .ZN(_03359_)
);

NAND2_X1 _08755_ (
  .A1(_03317_),
  .A2(\sresult[40][0] ),
  .ZN(_03360_)
);

NAND2_X1 _08756_ (
  .A1(_03359_),
  .A2(_03360_),
  .ZN(_00480_)
);

NAND2_X1 _08757_ (
  .A1(_03312_),
  .A2(\sresult[39][1] ),
  .ZN(_03361_)
);

NAND2_X1 _08758_ (
  .A1(_03355_),
  .A2(din_42[1]),
  .ZN(_03362_)
);

NAND2_X1 _08759_ (
  .A1(_03361_),
  .A2(_03362_),
  .ZN(_03363_)
);

NAND2_X1 _08760_ (
  .A1(_03363_),
  .A2(_03358_),
  .ZN(_03364_)
);

NAND2_X1 _08761_ (
  .A1(_03317_),
  .A2(\sresult[40][1] ),
  .ZN(_03365_)
);

NAND2_X1 _08762_ (
  .A1(_03364_),
  .A2(_03365_),
  .ZN(_00481_)
);

BUF_X4 _08763_ (
  .A(_03147_),
  .Z(_03366_)
);

NAND2_X1 _08764_ (
  .A1(_03366_),
  .A2(\sresult[39][2] ),
  .ZN(_03367_)
);

NAND2_X1 _08765_ (
  .A1(_03355_),
  .A2(din_42[2]),
  .ZN(_03368_)
);

NAND2_X1 _08766_ (
  .A1(_03367_),
  .A2(_03368_),
  .ZN(_03369_)
);

NAND2_X1 _08767_ (
  .A1(_03369_),
  .A2(_03358_),
  .ZN(_03370_)
);

BUF_X1 _08768_ (
  .A(_03208_),
  .Z(_03371_)
);

NAND2_X1 _08769_ (
  .A1(_03371_),
  .A2(\sresult[40][2] ),
  .ZN(_03372_)
);

NAND2_X1 _08770_ (
  .A1(_03370_),
  .A2(_03372_),
  .ZN(_00482_)
);

NAND2_X1 _08771_ (
  .A1(_03366_),
  .A2(\sresult[39][3] ),
  .ZN(_03373_)
);

NAND2_X1 _08772_ (
  .A1(_03355_),
  .A2(din_42[3]),
  .ZN(_03374_)
);

NAND2_X1 _08773_ (
  .A1(_03373_),
  .A2(_03374_),
  .ZN(_03375_)
);

NAND2_X1 _08774_ (
  .A1(_03375_),
  .A2(_03358_),
  .ZN(_03376_)
);

NAND2_X1 _08775_ (
  .A1(_03371_),
  .A2(\sresult[40][3] ),
  .ZN(_03377_)
);

NAND2_X1 _08776_ (
  .A1(_03376_),
  .A2(_03377_),
  .ZN(_00483_)
);

NAND2_X1 _08777_ (
  .A1(_03366_),
  .A2(\sresult[39][4] ),
  .ZN(_03378_)
);

NAND2_X1 _08778_ (
  .A1(_03355_),
  .A2(din_42[4]),
  .ZN(_03379_)
);

NAND2_X1 _08779_ (
  .A1(_03378_),
  .A2(_03379_),
  .ZN(_03380_)
);

NAND2_X1 _08780_ (
  .A1(_03380_),
  .A2(_03358_),
  .ZN(_03381_)
);

NAND2_X1 _08781_ (
  .A1(_03371_),
  .A2(\sresult[40][4] ),
  .ZN(_03382_)
);

NAND2_X1 _08782_ (
  .A1(_03381_),
  .A2(_03382_),
  .ZN(_00484_)
);

NAND2_X1 _08783_ (
  .A1(_03366_),
  .A2(\sresult[39][5] ),
  .ZN(_03383_)
);

NAND2_X1 _08784_ (
  .A1(_03355_),
  .A2(din_42[5]),
  .ZN(_03384_)
);

NAND2_X1 _08785_ (
  .A1(_03383_),
  .A2(_03384_),
  .ZN(_03385_)
);

NAND2_X1 _08786_ (
  .A1(_03385_),
  .A2(_03358_),
  .ZN(_03386_)
);

NAND2_X1 _08787_ (
  .A1(_03371_),
  .A2(\sresult[40][5] ),
  .ZN(_03387_)
);

NAND2_X1 _08788_ (
  .A1(_03386_),
  .A2(_03387_),
  .ZN(_00485_)
);

NAND2_X1 _08789_ (
  .A1(_03366_),
  .A2(\sresult[39][6] ),
  .ZN(_03388_)
);

NAND2_X1 _08790_ (
  .A1(_03355_),
  .A2(din_42[6]),
  .ZN(_03389_)
);

NAND2_X1 _08791_ (
  .A1(_03388_),
  .A2(_03389_),
  .ZN(_03390_)
);

NAND2_X1 _08792_ (
  .A1(_03390_),
  .A2(_03358_),
  .ZN(_03391_)
);

NAND2_X1 _08793_ (
  .A1(_03371_),
  .A2(\sresult[40][6] ),
  .ZN(_03392_)
);

NAND2_X1 _08794_ (
  .A1(_03391_),
  .A2(_03392_),
  .ZN(_00486_)
);

NAND2_X1 _08795_ (
  .A1(_03366_),
  .A2(\sresult[39][7] ),
  .ZN(_03393_)
);

NAND2_X1 _08796_ (
  .A1(_03355_),
  .A2(din_42[7]),
  .ZN(_03394_)
);

NAND2_X1 _08797_ (
  .A1(_03393_),
  .A2(_03394_),
  .ZN(_03395_)
);

NAND2_X1 _08798_ (
  .A1(_03395_),
  .A2(_03358_),
  .ZN(_03396_)
);

NAND2_X1 _08799_ (
  .A1(_03371_),
  .A2(\sresult[40][7] ),
  .ZN(_03397_)
);

NAND2_X1 _08800_ (
  .A1(_03396_),
  .A2(_03397_),
  .ZN(_00487_)
);

NAND2_X1 _08801_ (
  .A1(_03366_),
  .A2(\sresult[39][8] ),
  .ZN(_03398_)
);

NAND2_X1 _08802_ (
  .A1(_03355_),
  .A2(din_42[8]),
  .ZN(_03399_)
);

NAND2_X1 _08803_ (
  .A1(_03398_),
  .A2(_03399_),
  .ZN(_03400_)
);

NAND2_X1 _08804_ (
  .A1(_03400_),
  .A2(_03358_),
  .ZN(_03401_)
);

NAND2_X1 _08805_ (
  .A1(_03371_),
  .A2(\sresult[40][8] ),
  .ZN(_03402_)
);

NAND2_X1 _08806_ (
  .A1(_03401_),
  .A2(_03402_),
  .ZN(_00488_)
);

NAND2_X1 _08807_ (
  .A1(_03366_),
  .A2(\sresult[39][9] ),
  .ZN(_03403_)
);

NAND2_X1 _08808_ (
  .A1(_03355_),
  .A2(din_42[9]),
  .ZN(_03404_)
);

NAND2_X1 _08809_ (
  .A1(_03403_),
  .A2(_03404_),
  .ZN(_03405_)
);

NAND2_X1 _08810_ (
  .A1(_03405_),
  .A2(_03358_),
  .ZN(_03406_)
);

NAND2_X1 _08811_ (
  .A1(_03371_),
  .A2(\sresult[40][9] ),
  .ZN(_03407_)
);

NAND2_X1 _08812_ (
  .A1(_03406_),
  .A2(_03407_),
  .ZN(_00489_)
);

NAND2_X1 _08813_ (
  .A1(_03366_),
  .A2(\sresult[39][10] ),
  .ZN(_03408_)
);

BUF_X4 _08814_ (
  .A(_03191_),
  .Z(_03409_)
);

NAND2_X1 _08815_ (
  .A1(_03409_),
  .A2(din_42[10]),
  .ZN(_03410_)
);

NAND2_X1 _08816_ (
  .A1(_03408_),
  .A2(_03410_),
  .ZN(_03411_)
);

BUF_X2 _08817_ (
  .A(_03084_),
  .Z(_03412_)
);

NAND2_X1 _08818_ (
  .A1(_03411_),
  .A2(_03412_),
  .ZN(_03413_)
);

NAND2_X1 _08819_ (
  .A1(_03371_),
  .A2(\sresult[40][10] ),
  .ZN(_03414_)
);

NAND2_X1 _08820_ (
  .A1(_03413_),
  .A2(_03414_),
  .ZN(_00490_)
);

NAND2_X1 _08821_ (
  .A1(_03366_),
  .A2(\sresult[39][11] ),
  .ZN(_03415_)
);

NAND2_X1 _08822_ (
  .A1(_03409_),
  .A2(din_42[11]),
  .ZN(_03416_)
);

NAND2_X1 _08823_ (
  .A1(_03415_),
  .A2(_03416_),
  .ZN(_03417_)
);

NAND2_X1 _08824_ (
  .A1(_03417_),
  .A2(_03412_),
  .ZN(_03418_)
);

NAND2_X1 _08825_ (
  .A1(_03371_),
  .A2(\sresult[40][11] ),
  .ZN(_03419_)
);

NAND2_X1 _08826_ (
  .A1(_03418_),
  .A2(_03419_),
  .ZN(_00491_)
);

BUF_X4 _08827_ (
  .A(_03147_),
  .Z(_03420_)
);

NAND2_X1 _08828_ (
  .A1(_03420_),
  .A2(\sresult[40][0] ),
  .ZN(_03421_)
);

NAND2_X1 _08829_ (
  .A1(_03409_),
  .A2(din_51[0]),
  .ZN(_03422_)
);

NAND2_X1 _08830_ (
  .A1(_03421_),
  .A2(_03422_),
  .ZN(_03423_)
);

NAND2_X1 _08831_ (
  .A1(_03423_),
  .A2(_03412_),
  .ZN(_03424_)
);

BUF_X1 _08832_ (
  .A(_03208_),
  .Z(_03425_)
);

NAND2_X1 _08833_ (
  .A1(_03425_),
  .A2(\sresult[41][0] ),
  .ZN(_03426_)
);

NAND2_X1 _08834_ (
  .A1(_03424_),
  .A2(_03426_),
  .ZN(_00492_)
);

NAND2_X1 _08835_ (
  .A1(_03420_),
  .A2(\sresult[40][1] ),
  .ZN(_03427_)
);

NAND2_X1 _08836_ (
  .A1(_03409_),
  .A2(din_51[1]),
  .ZN(_03428_)
);

NAND2_X1 _08837_ (
  .A1(_03427_),
  .A2(_03428_),
  .ZN(_03429_)
);

NAND2_X1 _08838_ (
  .A1(_03429_),
  .A2(_03412_),
  .ZN(_03430_)
);

NAND2_X1 _08839_ (
  .A1(_03425_),
  .A2(\sresult[41][1] ),
  .ZN(_03431_)
);

NAND2_X1 _08840_ (
  .A1(_03430_),
  .A2(_03431_),
  .ZN(_00493_)
);

NAND2_X1 _08841_ (
  .A1(_03420_),
  .A2(\sresult[40][2] ),
  .ZN(_03432_)
);

NAND2_X1 _08842_ (
  .A1(_03409_),
  .A2(din_51[2]),
  .ZN(_03433_)
);

NAND2_X1 _08843_ (
  .A1(_03432_),
  .A2(_03433_),
  .ZN(_03434_)
);

NAND2_X1 _08844_ (
  .A1(_03434_),
  .A2(_03412_),
  .ZN(_03435_)
);

NAND2_X1 _08845_ (
  .A1(_03425_),
  .A2(\sresult[41][2] ),
  .ZN(_03436_)
);

NAND2_X1 _08846_ (
  .A1(_03435_),
  .A2(_03436_),
  .ZN(_00494_)
);

NAND2_X1 _08847_ (
  .A1(_03420_),
  .A2(\sresult[40][3] ),
  .ZN(_03437_)
);

NAND2_X1 _08848_ (
  .A1(_03409_),
  .A2(din_51[3]),
  .ZN(_03438_)
);

NAND2_X1 _08849_ (
  .A1(_03437_),
  .A2(_03438_),
  .ZN(_03439_)
);

NAND2_X1 _08850_ (
  .A1(_03439_),
  .A2(_03412_),
  .ZN(_03440_)
);

NAND2_X1 _08851_ (
  .A1(_03425_),
  .A2(\sresult[41][3] ),
  .ZN(_03441_)
);

NAND2_X1 _08852_ (
  .A1(_03440_),
  .A2(_03441_),
  .ZN(_00495_)
);

NAND2_X1 _08853_ (
  .A1(_03420_),
  .A2(\sresult[40][4] ),
  .ZN(_03442_)
);

NAND2_X1 _08854_ (
  .A1(_03409_),
  .A2(din_51[4]),
  .ZN(_03443_)
);

NAND2_X1 _08855_ (
  .A1(_03442_),
  .A2(_03443_),
  .ZN(_03444_)
);

NAND2_X1 _08856_ (
  .A1(_03444_),
  .A2(_03412_),
  .ZN(_03445_)
);

NAND2_X1 _08857_ (
  .A1(_03425_),
  .A2(\sresult[41][4] ),
  .ZN(_03446_)
);

NAND2_X1 _08858_ (
  .A1(_03445_),
  .A2(_03446_),
  .ZN(_00496_)
);

NAND2_X1 _08859_ (
  .A1(_03420_),
  .A2(\sresult[40][5] ),
  .ZN(_03447_)
);

NAND2_X1 _08860_ (
  .A1(_03409_),
  .A2(din_51[5]),
  .ZN(_03448_)
);

NAND2_X1 _08861_ (
  .A1(_03447_),
  .A2(_03448_),
  .ZN(_03449_)
);

NAND2_X1 _08862_ (
  .A1(_03449_),
  .A2(_03412_),
  .ZN(_03450_)
);

NAND2_X1 _08863_ (
  .A1(_03425_),
  .A2(\sresult[41][5] ),
  .ZN(_03451_)
);

NAND2_X1 _08864_ (
  .A1(_03450_),
  .A2(_03451_),
  .ZN(_00497_)
);

NAND2_X1 _08865_ (
  .A1(_03420_),
  .A2(\sresult[40][6] ),
  .ZN(_03452_)
);

NAND2_X1 _08866_ (
  .A1(_03409_),
  .A2(din_51[6]),
  .ZN(_03453_)
);

NAND2_X1 _08867_ (
  .A1(_03452_),
  .A2(_03453_),
  .ZN(_03454_)
);

NAND2_X1 _08868_ (
  .A1(_03454_),
  .A2(_03412_),
  .ZN(_03455_)
);

NAND2_X1 _08869_ (
  .A1(_03425_),
  .A2(\sresult[41][6] ),
  .ZN(_03456_)
);

NAND2_X1 _08870_ (
  .A1(_03455_),
  .A2(_03456_),
  .ZN(_00498_)
);

NAND2_X1 _08871_ (
  .A1(_03420_),
  .A2(\sresult[40][7] ),
  .ZN(_03457_)
);

NAND2_X1 _08872_ (
  .A1(_03409_),
  .A2(din_51[7]),
  .ZN(_03458_)
);

NAND2_X1 _08873_ (
  .A1(_03457_),
  .A2(_03458_),
  .ZN(_03459_)
);

NAND2_X1 _08874_ (
  .A1(_03459_),
  .A2(_03412_),
  .ZN(_03460_)
);

NAND2_X1 _08875_ (
  .A1(_03425_),
  .A2(\sresult[41][7] ),
  .ZN(_03461_)
);

NAND2_X1 _08876_ (
  .A1(_03460_),
  .A2(_03461_),
  .ZN(_00499_)
);

NAND2_X1 _08877_ (
  .A1(_03420_),
  .A2(\sresult[40][8] ),
  .ZN(_03462_)
);

BUF_X4 _08878_ (
  .A(_03191_),
  .Z(_03463_)
);

NAND2_X1 _08879_ (
  .A1(_03463_),
  .A2(din_51[8]),
  .ZN(_03464_)
);

NAND2_X1 _08880_ (
  .A1(_03462_),
  .A2(_03464_),
  .ZN(_03465_)
);

BUF_X2 _08881_ (
  .A(_03084_),
  .Z(_03466_)
);

NAND2_X1 _08882_ (
  .A1(_03465_),
  .A2(_03466_),
  .ZN(_03467_)
);

NAND2_X1 _08883_ (
  .A1(_03425_),
  .A2(\sresult[41][8] ),
  .ZN(_03468_)
);

NAND2_X1 _08884_ (
  .A1(_03467_),
  .A2(_03468_),
  .ZN(_00500_)
);

NAND2_X1 _08885_ (
  .A1(_03420_),
  .A2(\sresult[40][9] ),
  .ZN(_03469_)
);

NAND2_X1 _08886_ (
  .A1(_03463_),
  .A2(din_51[9]),
  .ZN(_03470_)
);

NAND2_X1 _08887_ (
  .A1(_03469_),
  .A2(_03470_),
  .ZN(_03471_)
);

NAND2_X1 _08888_ (
  .A1(_03471_),
  .A2(_03466_),
  .ZN(_03472_)
);

NAND2_X1 _08889_ (
  .A1(_03425_),
  .A2(\sresult[41][9] ),
  .ZN(_03473_)
);

NAND2_X1 _08890_ (
  .A1(_03472_),
  .A2(_03473_),
  .ZN(_00501_)
);

BUF_X4 _08891_ (
  .A(_03147_),
  .Z(_03474_)
);

NAND2_X1 _08892_ (
  .A1(_03474_),
  .A2(\sresult[40][10] ),
  .ZN(_03475_)
);

NAND2_X1 _08893_ (
  .A1(_03463_),
  .A2(din_51[10]),
  .ZN(_03476_)
);

NAND2_X1 _08894_ (
  .A1(_03475_),
  .A2(_03476_),
  .ZN(_03477_)
);

NAND2_X1 _08895_ (
  .A1(_03477_),
  .A2(_03466_),
  .ZN(_03478_)
);

BUF_X1 _08896_ (
  .A(_03208_),
  .Z(_03479_)
);

NAND2_X1 _08897_ (
  .A1(_03479_),
  .A2(\sresult[41][10] ),
  .ZN(_03480_)
);

NAND2_X1 _08898_ (
  .A1(_03478_),
  .A2(_03480_),
  .ZN(_00502_)
);

NAND2_X1 _08899_ (
  .A1(_03474_),
  .A2(\sresult[40][11] ),
  .ZN(_03481_)
);

NAND2_X1 _08900_ (
  .A1(_03463_),
  .A2(din_51[11]),
  .ZN(_03482_)
);

NAND2_X1 _08901_ (
  .A1(_03481_),
  .A2(_03482_),
  .ZN(_03483_)
);

NAND2_X1 _08902_ (
  .A1(_03483_),
  .A2(_03466_),
  .ZN(_03484_)
);

NAND2_X1 _08903_ (
  .A1(_03479_),
  .A2(\sresult[41][11] ),
  .ZN(_03485_)
);

NAND2_X1 _08904_ (
  .A1(_03484_),
  .A2(_03485_),
  .ZN(_00503_)
);

NAND2_X1 _08905_ (
  .A1(_03474_),
  .A2(\sresult[41][0] ),
  .ZN(_03486_)
);

NAND2_X1 _08906_ (
  .A1(_03463_),
  .A2(din_60[0]),
  .ZN(_03487_)
);

NAND2_X1 _08907_ (
  .A1(_03486_),
  .A2(_03487_),
  .ZN(_03488_)
);

NAND2_X1 _08908_ (
  .A1(_03488_),
  .A2(_03466_),
  .ZN(_03489_)
);

NAND2_X1 _08909_ (
  .A1(_03479_),
  .A2(\sresult[42][0] ),
  .ZN(_03490_)
);

NAND2_X1 _08910_ (
  .A1(_03489_),
  .A2(_03490_),
  .ZN(_00504_)
);

NAND2_X1 _08911_ (
  .A1(_03474_),
  .A2(\sresult[41][1] ),
  .ZN(_03491_)
);

NAND2_X1 _08912_ (
  .A1(_03463_),
  .A2(din_60[1]),
  .ZN(_03492_)
);

NAND2_X1 _08913_ (
  .A1(_03491_),
  .A2(_03492_),
  .ZN(_03493_)
);

NAND2_X1 _08914_ (
  .A1(_03493_),
  .A2(_03466_),
  .ZN(_03494_)
);

NAND2_X1 _08915_ (
  .A1(_03479_),
  .A2(\sresult[42][1] ),
  .ZN(_03495_)
);

NAND2_X1 _08916_ (
  .A1(_03494_),
  .A2(_03495_),
  .ZN(_00505_)
);

NAND2_X1 _08917_ (
  .A1(_03474_),
  .A2(\sresult[41][2] ),
  .ZN(_03496_)
);

NAND2_X1 _08918_ (
  .A1(_03463_),
  .A2(din_60[2]),
  .ZN(_03497_)
);

NAND2_X1 _08919_ (
  .A1(_03496_),
  .A2(_03497_),
  .ZN(_03498_)
);

NAND2_X1 _08920_ (
  .A1(_03498_),
  .A2(_03466_),
  .ZN(_03499_)
);

NAND2_X1 _08921_ (
  .A1(_03479_),
  .A2(\sresult[42][2] ),
  .ZN(_03500_)
);

NAND2_X1 _08922_ (
  .A1(_03499_),
  .A2(_03500_),
  .ZN(_00506_)
);

NAND2_X1 _08923_ (
  .A1(_03474_),
  .A2(\sresult[41][3] ),
  .ZN(_03501_)
);

NAND2_X1 _08924_ (
  .A1(_03463_),
  .A2(din_60[3]),
  .ZN(_03502_)
);

NAND2_X1 _08925_ (
  .A1(_03501_),
  .A2(_03502_),
  .ZN(_03503_)
);

NAND2_X1 _08926_ (
  .A1(_03503_),
  .A2(_03466_),
  .ZN(_03504_)
);

NAND2_X1 _08927_ (
  .A1(_03479_),
  .A2(\sresult[42][3] ),
  .ZN(_03505_)
);

NAND2_X1 _08928_ (
  .A1(_03504_),
  .A2(_03505_),
  .ZN(_00507_)
);

NAND2_X1 _08929_ (
  .A1(_03474_),
  .A2(\sresult[41][4] ),
  .ZN(_03506_)
);

NAND2_X1 _08930_ (
  .A1(_03463_),
  .A2(din_60[4]),
  .ZN(_03507_)
);

NAND2_X1 _08931_ (
  .A1(_03506_),
  .A2(_03507_),
  .ZN(_03508_)
);

NAND2_X1 _08932_ (
  .A1(_03508_),
  .A2(_03466_),
  .ZN(_03509_)
);

NAND2_X1 _08933_ (
  .A1(_03479_),
  .A2(\sresult[42][4] ),
  .ZN(_03510_)
);

NAND2_X1 _08934_ (
  .A1(_03509_),
  .A2(_03510_),
  .ZN(_00508_)
);

NAND2_X1 _08935_ (
  .A1(_03474_),
  .A2(\sresult[41][5] ),
  .ZN(_03511_)
);

NAND2_X1 _08936_ (
  .A1(_03463_),
  .A2(din_60[5]),
  .ZN(_03512_)
);

NAND2_X1 _08937_ (
  .A1(_03511_),
  .A2(_03512_),
  .ZN(_03513_)
);

NAND2_X1 _08938_ (
  .A1(_03513_),
  .A2(_03466_),
  .ZN(_03514_)
);

NAND2_X1 _08939_ (
  .A1(_03479_),
  .A2(\sresult[42][5] ),
  .ZN(_03515_)
);

NAND2_X1 _08940_ (
  .A1(_03514_),
  .A2(_03515_),
  .ZN(_00509_)
);

NAND2_X1 _08941_ (
  .A1(_03474_),
  .A2(\sresult[41][6] ),
  .ZN(_03516_)
);

BUF_X4 _08942_ (
  .A(_03191_),
  .Z(_03517_)
);

NAND2_X1 _08943_ (
  .A1(_03517_),
  .A2(din_60[6]),
  .ZN(_03518_)
);

NAND2_X1 _08944_ (
  .A1(_03516_),
  .A2(_03518_),
  .ZN(_03519_)
);

BUF_X2 _08945_ (
  .A(_03084_),
  .Z(_03520_)
);

NAND2_X1 _08946_ (
  .A1(_03519_),
  .A2(_03520_),
  .ZN(_03521_)
);

NAND2_X1 _08947_ (
  .A1(_03479_),
  .A2(\sresult[42][6] ),
  .ZN(_03522_)
);

NAND2_X1 _08948_ (
  .A1(_03521_),
  .A2(_03522_),
  .ZN(_00510_)
);

NAND2_X1 _08949_ (
  .A1(_03474_),
  .A2(\sresult[41][7] ),
  .ZN(_03523_)
);

NAND2_X1 _08950_ (
  .A1(_03517_),
  .A2(din_60[7]),
  .ZN(_03524_)
);

NAND2_X1 _08951_ (
  .A1(_03523_),
  .A2(_03524_),
  .ZN(_03525_)
);

NAND2_X1 _08952_ (
  .A1(_03525_),
  .A2(_03520_),
  .ZN(_03526_)
);

NAND2_X1 _08953_ (
  .A1(_03479_),
  .A2(\sresult[42][7] ),
  .ZN(_03527_)
);

NAND2_X1 _08954_ (
  .A1(_03526_),
  .A2(_03527_),
  .ZN(_00511_)
);

BUF_X4 _08955_ (
  .A(_03147_),
  .Z(_03528_)
);

NAND2_X1 _08956_ (
  .A1(_03528_),
  .A2(\sresult[41][8] ),
  .ZN(_03529_)
);

NAND2_X1 _08957_ (
  .A1(_03517_),
  .A2(din_60[8]),
  .ZN(_03530_)
);

NAND2_X1 _08958_ (
  .A1(_03529_),
  .A2(_03530_),
  .ZN(_03531_)
);

NAND2_X1 _08959_ (
  .A1(_03531_),
  .A2(_03520_),
  .ZN(_03532_)
);

BUF_X1 _08960_ (
  .A(_03208_),
  .Z(_03533_)
);

NAND2_X1 _08961_ (
  .A1(_03533_),
  .A2(\sresult[42][8] ),
  .ZN(_03534_)
);

NAND2_X1 _08962_ (
  .A1(_03532_),
  .A2(_03534_),
  .ZN(_00512_)
);

NAND2_X1 _08963_ (
  .A1(_03528_),
  .A2(\sresult[41][9] ),
  .ZN(_03535_)
);

NAND2_X1 _08964_ (
  .A1(_03517_),
  .A2(din_60[9]),
  .ZN(_03536_)
);

NAND2_X1 _08965_ (
  .A1(_03535_),
  .A2(_03536_),
  .ZN(_03537_)
);

NAND2_X1 _08966_ (
  .A1(_03537_),
  .A2(_03520_),
  .ZN(_03538_)
);

NAND2_X1 _08967_ (
  .A1(_03533_),
  .A2(\sresult[42][9] ),
  .ZN(_03539_)
);

NAND2_X1 _08968_ (
  .A1(_03538_),
  .A2(_03539_),
  .ZN(_00513_)
);

NAND2_X1 _08969_ (
  .A1(_03528_),
  .A2(\sresult[41][10] ),
  .ZN(_03540_)
);

NAND2_X1 _08970_ (
  .A1(_03517_),
  .A2(din_60[10]),
  .ZN(_03541_)
);

NAND2_X1 _08971_ (
  .A1(_03540_),
  .A2(_03541_),
  .ZN(_03542_)
);

NAND2_X1 _08972_ (
  .A1(_03542_),
  .A2(_03520_),
  .ZN(_03543_)
);

NAND2_X1 _08973_ (
  .A1(_03533_),
  .A2(\sresult[42][10] ),
  .ZN(_03544_)
);

NAND2_X1 _08974_ (
  .A1(_03543_),
  .A2(_03544_),
  .ZN(_00514_)
);

NAND2_X1 _08975_ (
  .A1(_03528_),
  .A2(\sresult[41][11] ),
  .ZN(_03545_)
);

NAND2_X1 _08976_ (
  .A1(_03517_),
  .A2(din_60[11]),
  .ZN(_03546_)
);

NAND2_X1 _08977_ (
  .A1(_03545_),
  .A2(_03546_),
  .ZN(_03547_)
);

NAND2_X1 _08978_ (
  .A1(_03547_),
  .A2(_03520_),
  .ZN(_03548_)
);

NAND2_X1 _08979_ (
  .A1(_03533_),
  .A2(\sresult[42][11] ),
  .ZN(_03549_)
);

NAND2_X1 _08980_ (
  .A1(_03548_),
  .A2(_03549_),
  .ZN(_00515_)
);

NAND2_X1 _08981_ (
  .A1(_03528_),
  .A2(\sresult[42][0] ),
  .ZN(_03550_)
);

NAND2_X1 _08982_ (
  .A1(_03517_),
  .A2(din_50[0]),
  .ZN(_03551_)
);

NAND2_X1 _08983_ (
  .A1(_03550_),
  .A2(_03551_),
  .ZN(_03552_)
);

NAND2_X1 _08984_ (
  .A1(_03552_),
  .A2(_03520_),
  .ZN(_03553_)
);

NAND2_X1 _08985_ (
  .A1(_03533_),
  .A2(\sresult[43][0] ),
  .ZN(_03554_)
);

NAND2_X1 _08986_ (
  .A1(_03553_),
  .A2(_03554_),
  .ZN(_00516_)
);

NAND2_X1 _08987_ (
  .A1(_03528_),
  .A2(\sresult[42][1] ),
  .ZN(_03555_)
);

NAND2_X1 _08988_ (
  .A1(_03517_),
  .A2(din_50[1]),
  .ZN(_03556_)
);

NAND2_X1 _08989_ (
  .A1(_03555_),
  .A2(_03556_),
  .ZN(_03557_)
);

NAND2_X1 _08990_ (
  .A1(_03557_),
  .A2(_03520_),
  .ZN(_03558_)
);

NAND2_X1 _08991_ (
  .A1(_03533_),
  .A2(\sresult[43][1] ),
  .ZN(_03559_)
);

NAND2_X1 _08992_ (
  .A1(_03558_),
  .A2(_03559_),
  .ZN(_00517_)
);

NAND2_X1 _08993_ (
  .A1(_03528_),
  .A2(\sresult[42][2] ),
  .ZN(_03560_)
);

NAND2_X1 _08994_ (
  .A1(_03517_),
  .A2(din_50[2]),
  .ZN(_03561_)
);

NAND2_X1 _08995_ (
  .A1(_03560_),
  .A2(_03561_),
  .ZN(_03562_)
);

NAND2_X1 _08996_ (
  .A1(_03562_),
  .A2(_03520_),
  .ZN(_03563_)
);

NAND2_X1 _08997_ (
  .A1(_03533_),
  .A2(\sresult[43][2] ),
  .ZN(_03564_)
);

NAND2_X1 _08998_ (
  .A1(_03563_),
  .A2(_03564_),
  .ZN(_00518_)
);

NAND2_X1 _08999_ (
  .A1(_03528_),
  .A2(\sresult[42][3] ),
  .ZN(_03565_)
);

NAND2_X1 _09000_ (
  .A1(_03517_),
  .A2(din_50[3]),
  .ZN(_03566_)
);

NAND2_X1 _09001_ (
  .A1(_03565_),
  .A2(_03566_),
  .ZN(_03567_)
);

NAND2_X1 _09002_ (
  .A1(_03567_),
  .A2(_03520_),
  .ZN(_03568_)
);

NAND2_X1 _09003_ (
  .A1(_03533_),
  .A2(\sresult[43][3] ),
  .ZN(_03569_)
);

NAND2_X1 _09004_ (
  .A1(_03568_),
  .A2(_03569_),
  .ZN(_00519_)
);

NAND2_X1 _09005_ (
  .A1(_03528_),
  .A2(\sresult[42][4] ),
  .ZN(_03570_)
);

BUF_X4 _09006_ (
  .A(_03191_),
  .Z(_03571_)
);

NAND2_X1 _09007_ (
  .A1(_03571_),
  .A2(din_50[4]),
  .ZN(_03572_)
);

NAND2_X1 _09008_ (
  .A1(_03570_),
  .A2(_03572_),
  .ZN(_03573_)
);

BUF_X2 _09009_ (
  .A(_03084_),
  .Z(_03574_)
);

NAND2_X1 _09010_ (
  .A1(_03573_),
  .A2(_03574_),
  .ZN(_03575_)
);

NAND2_X1 _09011_ (
  .A1(_03533_),
  .A2(\sresult[43][4] ),
  .ZN(_03576_)
);

NAND2_X1 _09012_ (
  .A1(_03575_),
  .A2(_03576_),
  .ZN(_00520_)
);

NAND2_X1 _09013_ (
  .A1(_03528_),
  .A2(\sresult[42][5] ),
  .ZN(_03577_)
);

NAND2_X1 _09014_ (
  .A1(_03571_),
  .A2(din_50[5]),
  .ZN(_03578_)
);

NAND2_X1 _09015_ (
  .A1(_03577_),
  .A2(_03578_),
  .ZN(_03579_)
);

NAND2_X1 _09016_ (
  .A1(_03579_),
  .A2(_03574_),
  .ZN(_03580_)
);

NAND2_X1 _09017_ (
  .A1(_03533_),
  .A2(\sresult[43][5] ),
  .ZN(_03581_)
);

NAND2_X1 _09018_ (
  .A1(_03580_),
  .A2(_03581_),
  .ZN(_00521_)
);

BUF_X4 _09019_ (
  .A(_03147_),
  .Z(_03582_)
);

NAND2_X1 _09020_ (
  .A1(_03582_),
  .A2(\sresult[42][6] ),
  .ZN(_03583_)
);

NAND2_X1 _09021_ (
  .A1(_03571_),
  .A2(din_50[6]),
  .ZN(_03584_)
);

NAND2_X1 _09022_ (
  .A1(_03583_),
  .A2(_03584_),
  .ZN(_03585_)
);

NAND2_X1 _09023_ (
  .A1(_03585_),
  .A2(_03574_),
  .ZN(_03586_)
);

BUF_X1 _09024_ (
  .A(_03208_),
  .Z(_03587_)
);

NAND2_X1 _09025_ (
  .A1(_03587_),
  .A2(\sresult[43][6] ),
  .ZN(_03588_)
);

NAND2_X1 _09026_ (
  .A1(_03586_),
  .A2(_03588_),
  .ZN(_00522_)
);

NAND2_X1 _09027_ (
  .A1(_03582_),
  .A2(\sresult[42][7] ),
  .ZN(_03589_)
);

NAND2_X1 _09028_ (
  .A1(_03571_),
  .A2(din_50[7]),
  .ZN(_03590_)
);

NAND2_X1 _09029_ (
  .A1(_03589_),
  .A2(_03590_),
  .ZN(_03591_)
);

NAND2_X1 _09030_ (
  .A1(_03591_),
  .A2(_03574_),
  .ZN(_03592_)
);

NAND2_X1 _09031_ (
  .A1(_03587_),
  .A2(\sresult[43][7] ),
  .ZN(_03593_)
);

NAND2_X1 _09032_ (
  .A1(_03592_),
  .A2(_03593_),
  .ZN(_00523_)
);

NAND2_X1 _09033_ (
  .A1(_03582_),
  .A2(\sresult[42][8] ),
  .ZN(_03594_)
);

NAND2_X1 _09034_ (
  .A1(_03571_),
  .A2(din_50[8]),
  .ZN(_03595_)
);

NAND2_X1 _09035_ (
  .A1(_03594_),
  .A2(_03595_),
  .ZN(_03596_)
);

NAND2_X1 _09036_ (
  .A1(_03596_),
  .A2(_03574_),
  .ZN(_03597_)
);

NAND2_X1 _09037_ (
  .A1(_03587_),
  .A2(\sresult[43][8] ),
  .ZN(_03598_)
);

NAND2_X1 _09038_ (
  .A1(_03597_),
  .A2(_03598_),
  .ZN(_00524_)
);

NAND2_X1 _09039_ (
  .A1(_03582_),
  .A2(\sresult[42][9] ),
  .ZN(_03599_)
);

NAND2_X1 _09040_ (
  .A1(_03571_),
  .A2(din_50[9]),
  .ZN(_03600_)
);

NAND2_X1 _09041_ (
  .A1(_03599_),
  .A2(_03600_),
  .ZN(_03601_)
);

NAND2_X1 _09042_ (
  .A1(_03601_),
  .A2(_03574_),
  .ZN(_03602_)
);

NAND2_X1 _09043_ (
  .A1(_03587_),
  .A2(\sresult[43][9] ),
  .ZN(_03603_)
);

NAND2_X1 _09044_ (
  .A1(_03602_),
  .A2(_03603_),
  .ZN(_00525_)
);

NAND2_X1 _09045_ (
  .A1(_03582_),
  .A2(\sresult[42][10] ),
  .ZN(_03604_)
);

NAND2_X1 _09046_ (
  .A1(_03571_),
  .A2(din_50[10]),
  .ZN(_03605_)
);

NAND2_X1 _09047_ (
  .A1(_03604_),
  .A2(_03605_),
  .ZN(_03606_)
);

NAND2_X1 _09048_ (
  .A1(_03606_),
  .A2(_03574_),
  .ZN(_03607_)
);

NAND2_X1 _09049_ (
  .A1(_03587_),
  .A2(\sresult[43][10] ),
  .ZN(_03608_)
);

NAND2_X1 _09050_ (
  .A1(_03607_),
  .A2(_03608_),
  .ZN(_00526_)
);

NAND2_X1 _09051_ (
  .A1(_03582_),
  .A2(\sresult[42][11] ),
  .ZN(_03609_)
);

NAND2_X1 _09052_ (
  .A1(_03571_),
  .A2(din_50[11]),
  .ZN(_03610_)
);

NAND2_X1 _09053_ (
  .A1(_03609_),
  .A2(_03610_),
  .ZN(_03611_)
);

NAND2_X1 _09054_ (
  .A1(_03611_),
  .A2(_03574_),
  .ZN(_03612_)
);

NAND2_X1 _09055_ (
  .A1(_03587_),
  .A2(\sresult[43][11] ),
  .ZN(_03613_)
);

NAND2_X1 _09056_ (
  .A1(_03612_),
  .A2(_03613_),
  .ZN(_00527_)
);

NAND2_X1 _09057_ (
  .A1(_03582_),
  .A2(\sresult[43][0] ),
  .ZN(_03614_)
);

NAND2_X1 _09058_ (
  .A1(_03571_),
  .A2(din_41[0]),
  .ZN(_03615_)
);

NAND2_X1 _09059_ (
  .A1(_03614_),
  .A2(_03615_),
  .ZN(_03616_)
);

NAND2_X1 _09060_ (
  .A1(_03616_),
  .A2(_03574_),
  .ZN(_03617_)
);

NAND2_X1 _09061_ (
  .A1(_03587_),
  .A2(\sresult[44][0] ),
  .ZN(_03618_)
);

NAND2_X1 _09062_ (
  .A1(_03617_),
  .A2(_03618_),
  .ZN(_00528_)
);

NAND2_X1 _09063_ (
  .A1(_03582_),
  .A2(\sresult[43][1] ),
  .ZN(_03619_)
);

NAND2_X1 _09064_ (
  .A1(_03571_),
  .A2(din_41[1]),
  .ZN(_03620_)
);

NAND2_X1 _09065_ (
  .A1(_03619_),
  .A2(_03620_),
  .ZN(_03621_)
);

NAND2_X1 _09066_ (
  .A1(_03621_),
  .A2(_03574_),
  .ZN(_03622_)
);

NAND2_X1 _09067_ (
  .A1(_03587_),
  .A2(\sresult[44][1] ),
  .ZN(_03623_)
);

NAND2_X1 _09068_ (
  .A1(_03622_),
  .A2(_03623_),
  .ZN(_00529_)
);

NAND2_X1 _09069_ (
  .A1(_03582_),
  .A2(\sresult[43][2] ),
  .ZN(_03624_)
);

BUF_X4 _09070_ (
  .A(_03191_),
  .Z(_03625_)
);

NAND2_X1 _09071_ (
  .A1(_03625_),
  .A2(din_41[2]),
  .ZN(_03626_)
);

NAND2_X1 _09072_ (
  .A1(_03624_),
  .A2(_03626_),
  .ZN(_03627_)
);

BUF_X4 _09073_ (
  .A(_00911_),
  .Z(_03628_)
);

BUF_X2 _09074_ (
  .A(_03628_),
  .Z(_03629_)
);

NAND2_X1 _09075_ (
  .A1(_03627_),
  .A2(_03629_),
  .ZN(_03630_)
);

NAND2_X1 _09076_ (
  .A1(_03587_),
  .A2(\sresult[44][2] ),
  .ZN(_03631_)
);

NAND2_X1 _09077_ (
  .A1(_03630_),
  .A2(_03631_),
  .ZN(_00530_)
);

NAND2_X1 _09078_ (
  .A1(_03582_),
  .A2(\sresult[43][3] ),
  .ZN(_03632_)
);

NAND2_X1 _09079_ (
  .A1(_03625_),
  .A2(din_41[3]),
  .ZN(_03633_)
);

NAND2_X1 _09080_ (
  .A1(_03632_),
  .A2(_03633_),
  .ZN(_03634_)
);

NAND2_X1 _09081_ (
  .A1(_03634_),
  .A2(_03629_),
  .ZN(_03635_)
);

NAND2_X1 _09082_ (
  .A1(_03587_),
  .A2(\sresult[44][3] ),
  .ZN(_03636_)
);

NAND2_X1 _09083_ (
  .A1(_03635_),
  .A2(_03636_),
  .ZN(_00531_)
);

BUF_X4 _09084_ (
  .A(_03147_),
  .Z(_03637_)
);

NAND2_X1 _09085_ (
  .A1(_03637_),
  .A2(\sresult[43][4] ),
  .ZN(_03638_)
);

NAND2_X1 _09086_ (
  .A1(_03625_),
  .A2(din_41[4]),
  .ZN(_03639_)
);

NAND2_X1 _09087_ (
  .A1(_03638_),
  .A2(_03639_),
  .ZN(_03640_)
);

NAND2_X1 _09088_ (
  .A1(_03640_),
  .A2(_03629_),
  .ZN(_03641_)
);

BUF_X1 _09089_ (
  .A(_03208_),
  .Z(_03642_)
);

NAND2_X1 _09090_ (
  .A1(_03642_),
  .A2(\sresult[44][4] ),
  .ZN(_03643_)
);

NAND2_X1 _09091_ (
  .A1(_03641_),
  .A2(_03643_),
  .ZN(_00532_)
);

NAND2_X1 _09092_ (
  .A1(_03637_),
  .A2(\sresult[43][5] ),
  .ZN(_03644_)
);

NAND2_X1 _09093_ (
  .A1(_03625_),
  .A2(din_41[5]),
  .ZN(_03645_)
);

NAND2_X1 _09094_ (
  .A1(_03644_),
  .A2(_03645_),
  .ZN(_03646_)
);

NAND2_X1 _09095_ (
  .A1(_03646_),
  .A2(_03629_),
  .ZN(_03647_)
);

NAND2_X1 _09096_ (
  .A1(_03642_),
  .A2(\sresult[44][5] ),
  .ZN(_03648_)
);

NAND2_X1 _09097_ (
  .A1(_03647_),
  .A2(_03648_),
  .ZN(_00533_)
);

NAND2_X1 _09098_ (
  .A1(_03637_),
  .A2(\sresult[43][6] ),
  .ZN(_03649_)
);

NAND2_X1 _09099_ (
  .A1(_03625_),
  .A2(din_41[6]),
  .ZN(_03650_)
);

NAND2_X1 _09100_ (
  .A1(_03649_),
  .A2(_03650_),
  .ZN(_03651_)
);

NAND2_X1 _09101_ (
  .A1(_03651_),
  .A2(_03629_),
  .ZN(_03652_)
);

NAND2_X1 _09102_ (
  .A1(_03642_),
  .A2(\sresult[44][6] ),
  .ZN(_03653_)
);

NAND2_X1 _09103_ (
  .A1(_03652_),
  .A2(_03653_),
  .ZN(_00534_)
);

NAND2_X1 _09104_ (
  .A1(_03637_),
  .A2(\sresult[43][7] ),
  .ZN(_03654_)
);

NAND2_X1 _09105_ (
  .A1(_03625_),
  .A2(din_41[7]),
  .ZN(_03655_)
);

NAND2_X1 _09106_ (
  .A1(_03654_),
  .A2(_03655_),
  .ZN(_03656_)
);

NAND2_X1 _09107_ (
  .A1(_03656_),
  .A2(_03629_),
  .ZN(_03657_)
);

NAND2_X1 _09108_ (
  .A1(_03642_),
  .A2(\sresult[44][7] ),
  .ZN(_03658_)
);

NAND2_X1 _09109_ (
  .A1(_03657_),
  .A2(_03658_),
  .ZN(_00535_)
);

NAND2_X1 _09110_ (
  .A1(_03637_),
  .A2(\sresult[43][8] ),
  .ZN(_03659_)
);

NAND2_X1 _09111_ (
  .A1(_03625_),
  .A2(din_41[8]),
  .ZN(_03660_)
);

NAND2_X1 _09112_ (
  .A1(_03659_),
  .A2(_03660_),
  .ZN(_03661_)
);

NAND2_X1 _09113_ (
  .A1(_03661_),
  .A2(_03629_),
  .ZN(_03662_)
);

NAND2_X1 _09114_ (
  .A1(_03642_),
  .A2(\sresult[44][8] ),
  .ZN(_03663_)
);

NAND2_X1 _09115_ (
  .A1(_03662_),
  .A2(_03663_),
  .ZN(_00536_)
);

NAND2_X1 _09116_ (
  .A1(_03637_),
  .A2(\sresult[43][9] ),
  .ZN(_03664_)
);

NAND2_X1 _09117_ (
  .A1(_03625_),
  .A2(din_41[9]),
  .ZN(_03665_)
);

NAND2_X1 _09118_ (
  .A1(_03664_),
  .A2(_03665_),
  .ZN(_03666_)
);

NAND2_X1 _09119_ (
  .A1(_03666_),
  .A2(_03629_),
  .ZN(_03667_)
);

NAND2_X1 _09120_ (
  .A1(_03642_),
  .A2(\sresult[44][9] ),
  .ZN(_03668_)
);

NAND2_X1 _09121_ (
  .A1(_03667_),
  .A2(_03668_),
  .ZN(_00537_)
);

NAND2_X1 _09122_ (
  .A1(_03637_),
  .A2(\sresult[43][10] ),
  .ZN(_03669_)
);

NAND2_X1 _09123_ (
  .A1(_03625_),
  .A2(din_41[10]),
  .ZN(_03670_)
);

NAND2_X1 _09124_ (
  .A1(_03669_),
  .A2(_03670_),
  .ZN(_03671_)
);

NAND2_X1 _09125_ (
  .A1(_03671_),
  .A2(_03629_),
  .ZN(_03672_)
);

NAND2_X1 _09126_ (
  .A1(_03642_),
  .A2(\sresult[44][10] ),
  .ZN(_03673_)
);

NAND2_X1 _09127_ (
  .A1(_03672_),
  .A2(_03673_),
  .ZN(_00538_)
);

NAND2_X1 _09128_ (
  .A1(_03637_),
  .A2(\sresult[43][11] ),
  .ZN(_03674_)
);

NAND2_X1 _09129_ (
  .A1(_03625_),
  .A2(din_41[11]),
  .ZN(_03675_)
);

NAND2_X1 _09130_ (
  .A1(_03674_),
  .A2(_03675_),
  .ZN(_03676_)
);

NAND2_X1 _09131_ (
  .A1(_03676_),
  .A2(_03629_),
  .ZN(_03677_)
);

NAND2_X1 _09132_ (
  .A1(_03642_),
  .A2(\sresult[44][11] ),
  .ZN(_03678_)
);

NAND2_X1 _09133_ (
  .A1(_03677_),
  .A2(_03678_),
  .ZN(_00539_)
);

NAND2_X1 _09134_ (
  .A1(_03637_),
  .A2(\sresult[44][0] ),
  .ZN(_03679_)
);

BUF_X4 _09135_ (
  .A(_03191_),
  .Z(_03680_)
);

NAND2_X1 _09136_ (
  .A1(_03680_),
  .A2(din_32[0]),
  .ZN(_03681_)
);

NAND2_X1 _09137_ (
  .A1(_03679_),
  .A2(_03681_),
  .ZN(_03682_)
);

BUF_X2 _09138_ (
  .A(_03628_),
  .Z(_03683_)
);

NAND2_X1 _09139_ (
  .A1(_03682_),
  .A2(_03683_),
  .ZN(_03684_)
);

NAND2_X1 _09140_ (
  .A1(_03642_),
  .A2(\sresult[45][0] ),
  .ZN(_03685_)
);

NAND2_X1 _09141_ (
  .A1(_03684_),
  .A2(_03685_),
  .ZN(_00540_)
);

NAND2_X1 _09142_ (
  .A1(_03637_),
  .A2(\sresult[44][1] ),
  .ZN(_03686_)
);

NAND2_X1 _09143_ (
  .A1(_03680_),
  .A2(din_32[1]),
  .ZN(_03687_)
);

NAND2_X1 _09144_ (
  .A1(_03686_),
  .A2(_03687_),
  .ZN(_03688_)
);

NAND2_X1 _09145_ (
  .A1(_03688_),
  .A2(_03683_),
  .ZN(_03689_)
);

NAND2_X1 _09146_ (
  .A1(_03642_),
  .A2(\sresult[45][1] ),
  .ZN(_03690_)
);

NAND2_X1 _09147_ (
  .A1(_03689_),
  .A2(_03690_),
  .ZN(_00541_)
);

BUF_X8 _09148_ (
  .A(_00799_),
  .Z(_03691_)
);

BUF_X4 _09149_ (
  .A(_03691_),
  .Z(_03692_)
);

NAND2_X1 _09150_ (
  .A1(_03692_),
  .A2(\sresult[44][2] ),
  .ZN(_03693_)
);

NAND2_X1 _09151_ (
  .A1(_03680_),
  .A2(din_32[2]),
  .ZN(_03694_)
);

NAND2_X1 _09152_ (
  .A1(_03693_),
  .A2(_03694_),
  .ZN(_03695_)
);

NAND2_X1 _09153_ (
  .A1(_03695_),
  .A2(_03683_),
  .ZN(_03696_)
);

BUF_X1 _09154_ (
  .A(_03208_),
  .Z(_03697_)
);

NAND2_X1 _09155_ (
  .A1(_03697_),
  .A2(\sresult[45][2] ),
  .ZN(_03698_)
);

NAND2_X1 _09156_ (
  .A1(_03696_),
  .A2(_03698_),
  .ZN(_00542_)
);

NAND2_X1 _09157_ (
  .A1(_03692_),
  .A2(\sresult[44][3] ),
  .ZN(_03699_)
);

NAND2_X1 _09158_ (
  .A1(_03680_),
  .A2(din_32[3]),
  .ZN(_03700_)
);

NAND2_X1 _09159_ (
  .A1(_03699_),
  .A2(_03700_),
  .ZN(_03701_)
);

NAND2_X1 _09160_ (
  .A1(_03701_),
  .A2(_03683_),
  .ZN(_03702_)
);

NAND2_X1 _09161_ (
  .A1(_03697_),
  .A2(\sresult[45][3] ),
  .ZN(_03703_)
);

NAND2_X1 _09162_ (
  .A1(_03702_),
  .A2(_03703_),
  .ZN(_00543_)
);

NAND2_X1 _09163_ (
  .A1(_03692_),
  .A2(\sresult[44][4] ),
  .ZN(_03704_)
);

NAND2_X1 _09164_ (
  .A1(_03680_),
  .A2(din_32[4]),
  .ZN(_03705_)
);

NAND2_X1 _09165_ (
  .A1(_03704_),
  .A2(_03705_),
  .ZN(_03706_)
);

NAND2_X1 _09166_ (
  .A1(_03706_),
  .A2(_03683_),
  .ZN(_03707_)
);

NAND2_X1 _09167_ (
  .A1(_03697_),
  .A2(\sresult[45][4] ),
  .ZN(_03708_)
);

NAND2_X1 _09168_ (
  .A1(_03707_),
  .A2(_03708_),
  .ZN(_00544_)
);

NAND2_X1 _09169_ (
  .A1(_03692_),
  .A2(\sresult[44][5] ),
  .ZN(_03709_)
);

NAND2_X1 _09170_ (
  .A1(_03680_),
  .A2(din_32[5]),
  .ZN(_03710_)
);

NAND2_X1 _09171_ (
  .A1(_03709_),
  .A2(_03710_),
  .ZN(_03711_)
);

NAND2_X1 _09172_ (
  .A1(_03711_),
  .A2(_03683_),
  .ZN(_03712_)
);

NAND2_X1 _09173_ (
  .A1(_03697_),
  .A2(\sresult[45][5] ),
  .ZN(_03713_)
);

NAND2_X1 _09174_ (
  .A1(_03712_),
  .A2(_03713_),
  .ZN(_00545_)
);

NAND2_X1 _09175_ (
  .A1(_03692_),
  .A2(\sresult[44][6] ),
  .ZN(_03714_)
);

NAND2_X1 _09176_ (
  .A1(_03680_),
  .A2(din_32[6]),
  .ZN(_03715_)
);

NAND2_X1 _09177_ (
  .A1(_03714_),
  .A2(_03715_),
  .ZN(_03716_)
);

NAND2_X1 _09178_ (
  .A1(_03716_),
  .A2(_03683_),
  .ZN(_03717_)
);

NAND2_X1 _09179_ (
  .A1(_03697_),
  .A2(\sresult[45][6] ),
  .ZN(_03718_)
);

NAND2_X1 _09180_ (
  .A1(_03717_),
  .A2(_03718_),
  .ZN(_00546_)
);

NAND2_X1 _09181_ (
  .A1(_03692_),
  .A2(\sresult[44][7] ),
  .ZN(_03719_)
);

NAND2_X1 _09182_ (
  .A1(_03680_),
  .A2(din_32[7]),
  .ZN(_03720_)
);

NAND2_X1 _09183_ (
  .A1(_03719_),
  .A2(_03720_),
  .ZN(_03721_)
);

NAND2_X1 _09184_ (
  .A1(_03721_),
  .A2(_03683_),
  .ZN(_03722_)
);

NAND2_X1 _09185_ (
  .A1(_03697_),
  .A2(\sresult[45][7] ),
  .ZN(_03723_)
);

NAND2_X1 _09186_ (
  .A1(_03722_),
  .A2(_03723_),
  .ZN(_00547_)
);

NAND2_X1 _09187_ (
  .A1(_03692_),
  .A2(\sresult[44][8] ),
  .ZN(_03724_)
);

NAND2_X1 _09188_ (
  .A1(_03680_),
  .A2(din_32[8]),
  .ZN(_03725_)
);

NAND2_X1 _09189_ (
  .A1(_03724_),
  .A2(_03725_),
  .ZN(_03726_)
);

NAND2_X1 _09190_ (
  .A1(_03726_),
  .A2(_03683_),
  .ZN(_03727_)
);

NAND2_X1 _09191_ (
  .A1(_03697_),
  .A2(\sresult[45][8] ),
  .ZN(_03728_)
);

NAND2_X1 _09192_ (
  .A1(_03727_),
  .A2(_03728_),
  .ZN(_00548_)
);

NAND2_X1 _09193_ (
  .A1(_03692_),
  .A2(\sresult[44][9] ),
  .ZN(_03729_)
);

NAND2_X1 _09194_ (
  .A1(_03680_),
  .A2(din_32[9]),
  .ZN(_03730_)
);

NAND2_X1 _09195_ (
  .A1(_03729_),
  .A2(_03730_),
  .ZN(_03731_)
);

NAND2_X1 _09196_ (
  .A1(_03731_),
  .A2(_03683_),
  .ZN(_03732_)
);

NAND2_X1 _09197_ (
  .A1(_03697_),
  .A2(\sresult[45][9] ),
  .ZN(_03733_)
);

NAND2_X1 _09198_ (
  .A1(_03732_),
  .A2(_03733_),
  .ZN(_00549_)
);

NAND2_X1 _09199_ (
  .A1(_03692_),
  .A2(\sresult[44][10] ),
  .ZN(_03734_)
);

BUF_X8 _09200_ (
  .A(_00770_),
  .Z(_03735_)
);

BUF_X4 _09201_ (
  .A(_03735_),
  .Z(_03736_)
);

NAND2_X1 _09202_ (
  .A1(_03736_),
  .A2(din_32[10]),
  .ZN(_03737_)
);

NAND2_X1 _09203_ (
  .A1(_03734_),
  .A2(_03737_),
  .ZN(_03738_)
);

BUF_X2 _09204_ (
  .A(_03628_),
  .Z(_03739_)
);

NAND2_X1 _09205_ (
  .A1(_03738_),
  .A2(_03739_),
  .ZN(_03740_)
);

NAND2_X1 _09206_ (
  .A1(_03697_),
  .A2(\sresult[45][10] ),
  .ZN(_03741_)
);

NAND2_X1 _09207_ (
  .A1(_03740_),
  .A2(_03741_),
  .ZN(_00550_)
);

NAND2_X1 _09208_ (
  .A1(_03692_),
  .A2(\sresult[44][11] ),
  .ZN(_03742_)
);

NAND2_X1 _09209_ (
  .A1(_03736_),
  .A2(din_32[11]),
  .ZN(_03743_)
);

NAND2_X1 _09210_ (
  .A1(_03742_),
  .A2(_03743_),
  .ZN(_03744_)
);

NAND2_X1 _09211_ (
  .A1(_03744_),
  .A2(_03739_),
  .ZN(_03745_)
);

NAND2_X1 _09212_ (
  .A1(_03697_),
  .A2(\sresult[45][11] ),
  .ZN(_03746_)
);

NAND2_X1 _09213_ (
  .A1(_03745_),
  .A2(_03746_),
  .ZN(_00551_)
);

BUF_X4 _09214_ (
  .A(_03691_),
  .Z(_03747_)
);

NAND2_X1 _09215_ (
  .A1(_03747_),
  .A2(\sresult[45][0] ),
  .ZN(_03748_)
);

NAND2_X1 _09216_ (
  .A1(_03736_),
  .A2(din_23[0]),
  .ZN(_03749_)
);

NAND2_X1 _09217_ (
  .A1(_03748_),
  .A2(_03749_),
  .ZN(_03750_)
);

NAND2_X1 _09218_ (
  .A1(_03750_),
  .A2(_03739_),
  .ZN(_03751_)
);

BUF_X8 _09219_ (
  .A(_00810_),
  .Z(_03752_)
);

BUF_X1 _09220_ (
  .A(_03752_),
  .Z(_03753_)
);

NAND2_X1 _09221_ (
  .A1(_03753_),
  .A2(\sresult[46][0] ),
  .ZN(_03754_)
);

NAND2_X1 _09222_ (
  .A1(_03751_),
  .A2(_03754_),
  .ZN(_00552_)
);

NAND2_X1 _09223_ (
  .A1(_03747_),
  .A2(\sresult[45][1] ),
  .ZN(_03755_)
);

NAND2_X1 _09224_ (
  .A1(_03736_),
  .A2(din_23[1]),
  .ZN(_03756_)
);

NAND2_X1 _09225_ (
  .A1(_03755_),
  .A2(_03756_),
  .ZN(_03757_)
);

NAND2_X1 _09226_ (
  .A1(_03757_),
  .A2(_03739_),
  .ZN(_03758_)
);

NAND2_X1 _09227_ (
  .A1(_03753_),
  .A2(\sresult[46][1] ),
  .ZN(_03759_)
);

NAND2_X1 _09228_ (
  .A1(_03758_),
  .A2(_03759_),
  .ZN(_00553_)
);

NAND2_X1 _09229_ (
  .A1(_03747_),
  .A2(\sresult[45][2] ),
  .ZN(_03760_)
);

NAND2_X1 _09230_ (
  .A1(_03736_),
  .A2(din_23[2]),
  .ZN(_03761_)
);

NAND2_X1 _09231_ (
  .A1(_03760_),
  .A2(_03761_),
  .ZN(_03762_)
);

NAND2_X1 _09232_ (
  .A1(_03762_),
  .A2(_03739_),
  .ZN(_03763_)
);

NAND2_X1 _09233_ (
  .A1(_03753_),
  .A2(\sresult[46][2] ),
  .ZN(_03764_)
);

NAND2_X1 _09234_ (
  .A1(_03763_),
  .A2(_03764_),
  .ZN(_00554_)
);

NAND2_X1 _09235_ (
  .A1(_03747_),
  .A2(\sresult[45][3] ),
  .ZN(_03765_)
);

NAND2_X1 _09236_ (
  .A1(_03736_),
  .A2(din_23[3]),
  .ZN(_03766_)
);

NAND2_X1 _09237_ (
  .A1(_03765_),
  .A2(_03766_),
  .ZN(_03767_)
);

NAND2_X1 _09238_ (
  .A1(_03767_),
  .A2(_03739_),
  .ZN(_03768_)
);

NAND2_X1 _09239_ (
  .A1(_03753_),
  .A2(\sresult[46][3] ),
  .ZN(_03769_)
);

NAND2_X1 _09240_ (
  .A1(_03768_),
  .A2(_03769_),
  .ZN(_00555_)
);

NAND2_X1 _09241_ (
  .A1(_03747_),
  .A2(\sresult[45][4] ),
  .ZN(_03770_)
);

NAND2_X1 _09242_ (
  .A1(_03736_),
  .A2(din_23[4]),
  .ZN(_03771_)
);

NAND2_X1 _09243_ (
  .A1(_03770_),
  .A2(_03771_),
  .ZN(_03772_)
);

NAND2_X1 _09244_ (
  .A1(_03772_),
  .A2(_03739_),
  .ZN(_03773_)
);

NAND2_X1 _09245_ (
  .A1(_03753_),
  .A2(\sresult[46][4] ),
  .ZN(_03774_)
);

NAND2_X1 _09246_ (
  .A1(_03773_),
  .A2(_03774_),
  .ZN(_00556_)
);

NAND2_X1 _09247_ (
  .A1(_03747_),
  .A2(\sresult[45][5] ),
  .ZN(_03775_)
);

NAND2_X1 _09248_ (
  .A1(_03736_),
  .A2(din_23[5]),
  .ZN(_03776_)
);

NAND2_X1 _09249_ (
  .A1(_03775_),
  .A2(_03776_),
  .ZN(_03777_)
);

NAND2_X1 _09250_ (
  .A1(_03777_),
  .A2(_03739_),
  .ZN(_03778_)
);

NAND2_X1 _09251_ (
  .A1(_03753_),
  .A2(\sresult[46][5] ),
  .ZN(_03779_)
);

NAND2_X1 _09252_ (
  .A1(_03778_),
  .A2(_03779_),
  .ZN(_00557_)
);

NAND2_X1 _09253_ (
  .A1(_03747_),
  .A2(\sresult[45][6] ),
  .ZN(_03780_)
);

NAND2_X1 _09254_ (
  .A1(_03736_),
  .A2(din_23[6]),
  .ZN(_03781_)
);

NAND2_X1 _09255_ (
  .A1(_03780_),
  .A2(_03781_),
  .ZN(_03782_)
);

NAND2_X1 _09256_ (
  .A1(_03782_),
  .A2(_03739_),
  .ZN(_03783_)
);

NAND2_X1 _09257_ (
  .A1(_03753_),
  .A2(\sresult[46][6] ),
  .ZN(_03784_)
);

NAND2_X1 _09258_ (
  .A1(_03783_),
  .A2(_03784_),
  .ZN(_00558_)
);

NAND2_X1 _09259_ (
  .A1(_03747_),
  .A2(\sresult[45][7] ),
  .ZN(_03785_)
);

NAND2_X1 _09260_ (
  .A1(_03736_),
  .A2(din_23[7]),
  .ZN(_03786_)
);

NAND2_X1 _09261_ (
  .A1(_03785_),
  .A2(_03786_),
  .ZN(_03787_)
);

NAND2_X1 _09262_ (
  .A1(_03787_),
  .A2(_03739_),
  .ZN(_03788_)
);

NAND2_X1 _09263_ (
  .A1(_03753_),
  .A2(\sresult[46][7] ),
  .ZN(_03789_)
);

NAND2_X1 _09264_ (
  .A1(_03788_),
  .A2(_03789_),
  .ZN(_00559_)
);

NAND2_X1 _09265_ (
  .A1(_03747_),
  .A2(\sresult[45][8] ),
  .ZN(_03790_)
);

BUF_X4 _09266_ (
  .A(_03735_),
  .Z(_03791_)
);

NAND2_X1 _09267_ (
  .A1(_03791_),
  .A2(din_23[8]),
  .ZN(_03792_)
);

NAND2_X1 _09268_ (
  .A1(_03790_),
  .A2(_03792_),
  .ZN(_03793_)
);

BUF_X2 _09269_ (
  .A(_03628_),
  .Z(_03794_)
);

NAND2_X1 _09270_ (
  .A1(_03793_),
  .A2(_03794_),
  .ZN(_03795_)
);

NAND2_X1 _09271_ (
  .A1(_03753_),
  .A2(\sresult[46][8] ),
  .ZN(_03796_)
);

NAND2_X1 _09272_ (
  .A1(_03795_),
  .A2(_03796_),
  .ZN(_00560_)
);

NAND2_X1 _09273_ (
  .A1(_03747_),
  .A2(\sresult[45][9] ),
  .ZN(_03797_)
);

NAND2_X1 _09274_ (
  .A1(_03791_),
  .A2(din_23[9]),
  .ZN(_03798_)
);

NAND2_X1 _09275_ (
  .A1(_03797_),
  .A2(_03798_),
  .ZN(_03799_)
);

NAND2_X1 _09276_ (
  .A1(_03799_),
  .A2(_03794_),
  .ZN(_03800_)
);

NAND2_X1 _09277_ (
  .A1(_03753_),
  .A2(\sresult[46][9] ),
  .ZN(_03801_)
);

NAND2_X1 _09278_ (
  .A1(_03800_),
  .A2(_03801_),
  .ZN(_00561_)
);

BUF_X4 _09279_ (
  .A(_03691_),
  .Z(_03802_)
);

NAND2_X1 _09280_ (
  .A1(_03802_),
  .A2(\sresult[45][10] ),
  .ZN(_03803_)
);

NAND2_X1 _09281_ (
  .A1(_03791_),
  .A2(din_23[10]),
  .ZN(_03804_)
);

NAND2_X1 _09282_ (
  .A1(_03803_),
  .A2(_03804_),
  .ZN(_03805_)
);

NAND2_X1 _09283_ (
  .A1(_03805_),
  .A2(_03794_),
  .ZN(_03806_)
);

BUF_X1 _09284_ (
  .A(_03752_),
  .Z(_03807_)
);

NAND2_X1 _09285_ (
  .A1(_03807_),
  .A2(\sresult[46][10] ),
  .ZN(_03808_)
);

NAND2_X1 _09286_ (
  .A1(_03806_),
  .A2(_03808_),
  .ZN(_00562_)
);

NAND2_X1 _09287_ (
  .A1(_03802_),
  .A2(\sresult[45][11] ),
  .ZN(_03809_)
);

NAND2_X1 _09288_ (
  .A1(_03791_),
  .A2(din_23[11]),
  .ZN(_03810_)
);

NAND2_X1 _09289_ (
  .A1(_03809_),
  .A2(_03810_),
  .ZN(_03811_)
);

NAND2_X1 _09290_ (
  .A1(_03811_),
  .A2(_03794_),
  .ZN(_03812_)
);

NAND2_X1 _09291_ (
  .A1(_03807_),
  .A2(\sresult[46][11] ),
  .ZN(_03813_)
);

NAND2_X1 _09292_ (
  .A1(_03812_),
  .A2(_03813_),
  .ZN(_00563_)
);

NAND2_X1 _09293_ (
  .A1(_03802_),
  .A2(\sresult[46][0] ),
  .ZN(_03814_)
);

NAND2_X1 _09294_ (
  .A1(_03791_),
  .A2(din_14[0]),
  .ZN(_03815_)
);

NAND2_X1 _09295_ (
  .A1(_03814_),
  .A2(_03815_),
  .ZN(_03816_)
);

NAND2_X1 _09296_ (
  .A1(_03816_),
  .A2(_03794_),
  .ZN(_03817_)
);

NAND2_X1 _09297_ (
  .A1(_03807_),
  .A2(\sresult[47][0] ),
  .ZN(_03818_)
);

NAND2_X1 _09298_ (
  .A1(_03817_),
  .A2(_03818_),
  .ZN(_00564_)
);

NAND2_X1 _09299_ (
  .A1(_03802_),
  .A2(\sresult[46][1] ),
  .ZN(_03819_)
);

NAND2_X1 _09300_ (
  .A1(_03791_),
  .A2(din_14[1]),
  .ZN(_03820_)
);

NAND2_X1 _09301_ (
  .A1(_03819_),
  .A2(_03820_),
  .ZN(_03821_)
);

NAND2_X1 _09302_ (
  .A1(_03821_),
  .A2(_03794_),
  .ZN(_03822_)
);

NAND2_X1 _09303_ (
  .A1(_03807_),
  .A2(\sresult[47][1] ),
  .ZN(_03823_)
);

NAND2_X1 _09304_ (
  .A1(_03822_),
  .A2(_03823_),
  .ZN(_00565_)
);

NAND2_X1 _09305_ (
  .A1(_03802_),
  .A2(\sresult[46][2] ),
  .ZN(_03824_)
);

NAND2_X1 _09306_ (
  .A1(_03791_),
  .A2(din_14[2]),
  .ZN(_03825_)
);

NAND2_X1 _09307_ (
  .A1(_03824_),
  .A2(_03825_),
  .ZN(_03826_)
);

NAND2_X1 _09308_ (
  .A1(_03826_),
  .A2(_03794_),
  .ZN(_03827_)
);

NAND2_X1 _09309_ (
  .A1(_03807_),
  .A2(\sresult[47][2] ),
  .ZN(_03828_)
);

NAND2_X1 _09310_ (
  .A1(_03827_),
  .A2(_03828_),
  .ZN(_00566_)
);

NAND2_X1 _09311_ (
  .A1(_03802_),
  .A2(\sresult[46][3] ),
  .ZN(_03829_)
);

NAND2_X1 _09312_ (
  .A1(_03791_),
  .A2(din_14[3]),
  .ZN(_03830_)
);

NAND2_X1 _09313_ (
  .A1(_03829_),
  .A2(_03830_),
  .ZN(_03831_)
);

NAND2_X1 _09314_ (
  .A1(_03831_),
  .A2(_03794_),
  .ZN(_03832_)
);

NAND2_X1 _09315_ (
  .A1(_03807_),
  .A2(\sresult[47][3] ),
  .ZN(_03833_)
);

NAND2_X1 _09316_ (
  .A1(_03832_),
  .A2(_03833_),
  .ZN(_00567_)
);

NAND2_X1 _09317_ (
  .A1(_03802_),
  .A2(\sresult[46][4] ),
  .ZN(_03834_)
);

NAND2_X1 _09318_ (
  .A1(_03791_),
  .A2(din_14[4]),
  .ZN(_03835_)
);

NAND2_X1 _09319_ (
  .A1(_03834_),
  .A2(_03835_),
  .ZN(_03836_)
);

NAND2_X1 _09320_ (
  .A1(_03836_),
  .A2(_03794_),
  .ZN(_03837_)
);

NAND2_X1 _09321_ (
  .A1(_03807_),
  .A2(\sresult[47][4] ),
  .ZN(_03838_)
);

NAND2_X1 _09322_ (
  .A1(_03837_),
  .A2(_03838_),
  .ZN(_00568_)
);

NAND2_X1 _09323_ (
  .A1(_03802_),
  .A2(\sresult[46][5] ),
  .ZN(_03839_)
);

NAND2_X1 _09324_ (
  .A1(_03791_),
  .A2(din_14[5]),
  .ZN(_03840_)
);

NAND2_X1 _09325_ (
  .A1(_03839_),
  .A2(_03840_),
  .ZN(_03841_)
);

NAND2_X1 _09326_ (
  .A1(_03841_),
  .A2(_03794_),
  .ZN(_03842_)
);

NAND2_X1 _09327_ (
  .A1(_03807_),
  .A2(\sresult[47][5] ),
  .ZN(_03843_)
);

NAND2_X1 _09328_ (
  .A1(_03842_),
  .A2(_03843_),
  .ZN(_00569_)
);

NAND2_X1 _09329_ (
  .A1(_03802_),
  .A2(\sresult[46][6] ),
  .ZN(_03844_)
);

BUF_X4 _09330_ (
  .A(_03735_),
  .Z(_03845_)
);

NAND2_X1 _09331_ (
  .A1(_03845_),
  .A2(din_14[6]),
  .ZN(_03846_)
);

NAND2_X1 _09332_ (
  .A1(_03844_),
  .A2(_03846_),
  .ZN(_03847_)
);

BUF_X2 _09333_ (
  .A(_03628_),
  .Z(_03848_)
);

NAND2_X1 _09334_ (
  .A1(_03847_),
  .A2(_03848_),
  .ZN(_03849_)
);

NAND2_X1 _09335_ (
  .A1(_03807_),
  .A2(\sresult[47][6] ),
  .ZN(_03850_)
);

NAND2_X1 _09336_ (
  .A1(_03849_),
  .A2(_03850_),
  .ZN(_00570_)
);

NAND2_X1 _09337_ (
  .A1(_03802_),
  .A2(\sresult[46][7] ),
  .ZN(_03851_)
);

NAND2_X1 _09338_ (
  .A1(_03845_),
  .A2(din_14[7]),
  .ZN(_03852_)
);

NAND2_X1 _09339_ (
  .A1(_03851_),
  .A2(_03852_),
  .ZN(_03853_)
);

NAND2_X1 _09340_ (
  .A1(_03853_),
  .A2(_03848_),
  .ZN(_03854_)
);

NAND2_X1 _09341_ (
  .A1(_03807_),
  .A2(\sresult[47][7] ),
  .ZN(_03855_)
);

NAND2_X1 _09342_ (
  .A1(_03854_),
  .A2(_03855_),
  .ZN(_00571_)
);

BUF_X4 _09343_ (
  .A(_03691_),
  .Z(_03856_)
);

NAND2_X1 _09344_ (
  .A1(_03856_),
  .A2(\sresult[46][8] ),
  .ZN(_03857_)
);

NAND2_X1 _09345_ (
  .A1(_03845_),
  .A2(din_14[8]),
  .ZN(_03858_)
);

NAND2_X1 _09346_ (
  .A1(_03857_),
  .A2(_03858_),
  .ZN(_03859_)
);

NAND2_X1 _09347_ (
  .A1(_03859_),
  .A2(_03848_),
  .ZN(_03860_)
);

BUF_X1 _09348_ (
  .A(_03752_),
  .Z(_03861_)
);

NAND2_X1 _09349_ (
  .A1(_03861_),
  .A2(\sresult[47][8] ),
  .ZN(_03862_)
);

NAND2_X1 _09350_ (
  .A1(_03860_),
  .A2(_03862_),
  .ZN(_00572_)
);

NAND2_X1 _09351_ (
  .A1(_03856_),
  .A2(\sresult[46][9] ),
  .ZN(_03863_)
);

NAND2_X1 _09352_ (
  .A1(_03845_),
  .A2(din_14[9]),
  .ZN(_03864_)
);

NAND2_X1 _09353_ (
  .A1(_03863_),
  .A2(_03864_),
  .ZN(_03865_)
);

NAND2_X1 _09354_ (
  .A1(_03865_),
  .A2(_03848_),
  .ZN(_03866_)
);

NAND2_X1 _09355_ (
  .A1(_03861_),
  .A2(\sresult[47][9] ),
  .ZN(_03867_)
);

NAND2_X1 _09356_ (
  .A1(_03866_),
  .A2(_03867_),
  .ZN(_00573_)
);

NAND2_X1 _09357_ (
  .A1(_03856_),
  .A2(\sresult[46][10] ),
  .ZN(_03868_)
);

NAND2_X1 _09358_ (
  .A1(_03845_),
  .A2(din_14[10]),
  .ZN(_03869_)
);

NAND2_X1 _09359_ (
  .A1(_03868_),
  .A2(_03869_),
  .ZN(_03870_)
);

NAND2_X1 _09360_ (
  .A1(_03870_),
  .A2(_03848_),
  .ZN(_03871_)
);

NAND2_X1 _09361_ (
  .A1(_03861_),
  .A2(\sresult[47][10] ),
  .ZN(_03872_)
);

NAND2_X1 _09362_ (
  .A1(_03871_),
  .A2(_03872_),
  .ZN(_00574_)
);

NAND2_X1 _09363_ (
  .A1(_03856_),
  .A2(\sresult[46][11] ),
  .ZN(_03873_)
);

NAND2_X1 _09364_ (
  .A1(_03845_),
  .A2(din_14[11]),
  .ZN(_03874_)
);

NAND2_X1 _09365_ (
  .A1(_03873_),
  .A2(_03874_),
  .ZN(_03875_)
);

NAND2_X1 _09366_ (
  .A1(_03875_),
  .A2(_03848_),
  .ZN(_03876_)
);

NAND2_X1 _09367_ (
  .A1(_03861_),
  .A2(\sresult[47][11] ),
  .ZN(_03877_)
);

NAND2_X1 _09368_ (
  .A1(_03876_),
  .A2(_03877_),
  .ZN(_00575_)
);

NAND2_X1 _09369_ (
  .A1(_03856_),
  .A2(\sresult[47][0] ),
  .ZN(_03878_)
);

NAND2_X1 _09370_ (
  .A1(_03845_),
  .A2(din_05[0]),
  .ZN(_03879_)
);

NAND2_X1 _09371_ (
  .A1(_03878_),
  .A2(_03879_),
  .ZN(_03880_)
);

NAND2_X1 _09372_ (
  .A1(_03880_),
  .A2(_03848_),
  .ZN(_03881_)
);

NAND2_X1 _09373_ (
  .A1(_03861_),
  .A2(\sresult[48][0] ),
  .ZN(_03882_)
);

NAND2_X1 _09374_ (
  .A1(_03881_),
  .A2(_03882_),
  .ZN(_00576_)
);

NAND2_X1 _09375_ (
  .A1(_03856_),
  .A2(\sresult[47][1] ),
  .ZN(_03883_)
);

NAND2_X1 _09376_ (
  .A1(_03845_),
  .A2(din_05[1]),
  .ZN(_03884_)
);

NAND2_X1 _09377_ (
  .A1(_03883_),
  .A2(_03884_),
  .ZN(_03885_)
);

NAND2_X1 _09378_ (
  .A1(_03885_),
  .A2(_03848_),
  .ZN(_03886_)
);

NAND2_X1 _09379_ (
  .A1(_03861_),
  .A2(\sresult[48][1] ),
  .ZN(_03887_)
);

NAND2_X1 _09380_ (
  .A1(_03886_),
  .A2(_03887_),
  .ZN(_00577_)
);

NAND2_X1 _09381_ (
  .A1(_03856_),
  .A2(\sresult[47][2] ),
  .ZN(_03888_)
);

NAND2_X1 _09382_ (
  .A1(_03845_),
  .A2(din_05[2]),
  .ZN(_03889_)
);

NAND2_X1 _09383_ (
  .A1(_03888_),
  .A2(_03889_),
  .ZN(_03890_)
);

NAND2_X1 _09384_ (
  .A1(_03890_),
  .A2(_03848_),
  .ZN(_03891_)
);

NAND2_X1 _09385_ (
  .A1(_03861_),
  .A2(\sresult[48][2] ),
  .ZN(_03892_)
);

NAND2_X1 _09386_ (
  .A1(_03891_),
  .A2(_03892_),
  .ZN(_00578_)
);

NAND2_X1 _09387_ (
  .A1(_03856_),
  .A2(\sresult[47][3] ),
  .ZN(_03893_)
);

NAND2_X1 _09388_ (
  .A1(_03845_),
  .A2(din_05[3]),
  .ZN(_03894_)
);

NAND2_X1 _09389_ (
  .A1(_03893_),
  .A2(_03894_),
  .ZN(_03895_)
);

NAND2_X1 _09390_ (
  .A1(_03895_),
  .A2(_03848_),
  .ZN(_03896_)
);

NAND2_X1 _09391_ (
  .A1(_03861_),
  .A2(\sresult[48][3] ),
  .ZN(_03897_)
);

NAND2_X1 _09392_ (
  .A1(_03896_),
  .A2(_03897_),
  .ZN(_00579_)
);

NAND2_X1 _09393_ (
  .A1(_03856_),
  .A2(\sresult[47][4] ),
  .ZN(_03898_)
);

BUF_X4 _09394_ (
  .A(_03735_),
  .Z(_03899_)
);

NAND2_X1 _09395_ (
  .A1(_03899_),
  .A2(din_05[4]),
  .ZN(_03900_)
);

NAND2_X1 _09396_ (
  .A1(_03898_),
  .A2(_03900_),
  .ZN(_03901_)
);

BUF_X2 _09397_ (
  .A(_03628_),
  .Z(_03902_)
);

NAND2_X1 _09398_ (
  .A1(_03901_),
  .A2(_03902_),
  .ZN(_03903_)
);

NAND2_X1 _09399_ (
  .A1(_03861_),
  .A2(\sresult[48][4] ),
  .ZN(_03904_)
);

NAND2_X1 _09400_ (
  .A1(_03903_),
  .A2(_03904_),
  .ZN(_00580_)
);

NAND2_X1 _09401_ (
  .A1(_03856_),
  .A2(\sresult[47][5] ),
  .ZN(_03905_)
);

NAND2_X1 _09402_ (
  .A1(_03899_),
  .A2(din_05[5]),
  .ZN(_03906_)
);

NAND2_X1 _09403_ (
  .A1(_03905_),
  .A2(_03906_),
  .ZN(_03907_)
);

NAND2_X1 _09404_ (
  .A1(_03907_),
  .A2(_03902_),
  .ZN(_03908_)
);

NAND2_X1 _09405_ (
  .A1(_03861_),
  .A2(\sresult[48][5] ),
  .ZN(_03909_)
);

NAND2_X1 _09406_ (
  .A1(_03908_),
  .A2(_03909_),
  .ZN(_00581_)
);

BUF_X4 _09407_ (
  .A(_03691_),
  .Z(_03910_)
);

NAND2_X1 _09408_ (
  .A1(_03910_),
  .A2(\sresult[47][6] ),
  .ZN(_03911_)
);

NAND2_X1 _09409_ (
  .A1(_03899_),
  .A2(din_05[6]),
  .ZN(_03912_)
);

NAND2_X1 _09410_ (
  .A1(_03911_),
  .A2(_03912_),
  .ZN(_03913_)
);

NAND2_X1 _09411_ (
  .A1(_03913_),
  .A2(_03902_),
  .ZN(_03914_)
);

BUF_X1 _09412_ (
  .A(_03752_),
  .Z(_03915_)
);

NAND2_X1 _09413_ (
  .A1(_03915_),
  .A2(\sresult[48][6] ),
  .ZN(_03916_)
);

NAND2_X1 _09414_ (
  .A1(_03914_),
  .A2(_03916_),
  .ZN(_00582_)
);

NAND2_X1 _09415_ (
  .A1(_03910_),
  .A2(\sresult[47][7] ),
  .ZN(_03917_)
);

NAND2_X1 _09416_ (
  .A1(_03899_),
  .A2(din_05[7]),
  .ZN(_03918_)
);

NAND2_X1 _09417_ (
  .A1(_03917_),
  .A2(_03918_),
  .ZN(_03919_)
);

NAND2_X1 _09418_ (
  .A1(_03919_),
  .A2(_03902_),
  .ZN(_03920_)
);

NAND2_X1 _09419_ (
  .A1(_03915_),
  .A2(\sresult[48][7] ),
  .ZN(_03921_)
);

NAND2_X1 _09420_ (
  .A1(_03920_),
  .A2(_03921_),
  .ZN(_00583_)
);

NAND2_X1 _09421_ (
  .A1(_03910_),
  .A2(\sresult[47][8] ),
  .ZN(_03922_)
);

NAND2_X1 _09422_ (
  .A1(_03899_),
  .A2(din_05[8]),
  .ZN(_03923_)
);

NAND2_X1 _09423_ (
  .A1(_03922_),
  .A2(_03923_),
  .ZN(_03924_)
);

NAND2_X1 _09424_ (
  .A1(_03924_),
  .A2(_03902_),
  .ZN(_03925_)
);

NAND2_X1 _09425_ (
  .A1(_03915_),
  .A2(\sresult[48][8] ),
  .ZN(_03926_)
);

NAND2_X1 _09426_ (
  .A1(_03925_),
  .A2(_03926_),
  .ZN(_00584_)
);

NAND2_X1 _09427_ (
  .A1(_03910_),
  .A2(\sresult[47][9] ),
  .ZN(_03927_)
);

NAND2_X1 _09428_ (
  .A1(_03899_),
  .A2(din_05[9]),
  .ZN(_03928_)
);

NAND2_X1 _09429_ (
  .A1(_03927_),
  .A2(_03928_),
  .ZN(_03929_)
);

NAND2_X1 _09430_ (
  .A1(_03929_),
  .A2(_03902_),
  .ZN(_03930_)
);

NAND2_X1 _09431_ (
  .A1(_03915_),
  .A2(\sresult[48][9] ),
  .ZN(_03931_)
);

NAND2_X1 _09432_ (
  .A1(_03930_),
  .A2(_03931_),
  .ZN(_00585_)
);

NAND2_X1 _09433_ (
  .A1(_03910_),
  .A2(\sresult[47][10] ),
  .ZN(_03932_)
);

NAND2_X1 _09434_ (
  .A1(_03899_),
  .A2(din_05[10]),
  .ZN(_03933_)
);

NAND2_X1 _09435_ (
  .A1(_03932_),
  .A2(_03933_),
  .ZN(_03934_)
);

NAND2_X1 _09436_ (
  .A1(_03934_),
  .A2(_03902_),
  .ZN(_03935_)
);

NAND2_X1 _09437_ (
  .A1(_03915_),
  .A2(\sresult[48][10] ),
  .ZN(_03936_)
);

NAND2_X1 _09438_ (
  .A1(_03935_),
  .A2(_03936_),
  .ZN(_00586_)
);

NAND2_X1 _09439_ (
  .A1(_03910_),
  .A2(\sresult[47][11] ),
  .ZN(_03937_)
);

NAND2_X1 _09440_ (
  .A1(_03899_),
  .A2(din_05[11]),
  .ZN(_03938_)
);

NAND2_X1 _09441_ (
  .A1(_03937_),
  .A2(_03938_),
  .ZN(_03939_)
);

NAND2_X1 _09442_ (
  .A1(_03939_),
  .A2(_03902_),
  .ZN(_03940_)
);

NAND2_X1 _09443_ (
  .A1(_03915_),
  .A2(\sresult[48][11] ),
  .ZN(_03941_)
);

NAND2_X1 _09444_ (
  .A1(_03940_),
  .A2(_03941_),
  .ZN(_00587_)
);

NAND2_X1 _09445_ (
  .A1(_03910_),
  .A2(\sresult[48][0] ),
  .ZN(_03942_)
);

NAND2_X1 _09446_ (
  .A1(_03899_),
  .A2(din_04[0]),
  .ZN(_03943_)
);

NAND2_X1 _09447_ (
  .A1(_03942_),
  .A2(_03943_),
  .ZN(_03944_)
);

NAND2_X1 _09448_ (
  .A1(_03944_),
  .A2(_03902_),
  .ZN(_03945_)
);

NAND2_X1 _09449_ (
  .A1(_03915_),
  .A2(\sresult[49][0] ),
  .ZN(_03946_)
);

NAND2_X1 _09450_ (
  .A1(_03945_),
  .A2(_03946_),
  .ZN(_00588_)
);

NAND2_X1 _09451_ (
  .A1(_03910_),
  .A2(\sresult[48][1] ),
  .ZN(_03947_)
);

NAND2_X1 _09452_ (
  .A1(_03899_),
  .A2(din_04[1]),
  .ZN(_03948_)
);

NAND2_X1 _09453_ (
  .A1(_03947_),
  .A2(_03948_),
  .ZN(_03949_)
);

NAND2_X1 _09454_ (
  .A1(_03949_),
  .A2(_03902_),
  .ZN(_03950_)
);

NAND2_X1 _09455_ (
  .A1(_03915_),
  .A2(\sresult[49][1] ),
  .ZN(_03951_)
);

NAND2_X1 _09456_ (
  .A1(_03950_),
  .A2(_03951_),
  .ZN(_00589_)
);

NAND2_X1 _09457_ (
  .A1(_03910_),
  .A2(\sresult[48][2] ),
  .ZN(_03952_)
);

BUF_X4 _09458_ (
  .A(_03735_),
  .Z(_03953_)
);

NAND2_X1 _09459_ (
  .A1(_03953_),
  .A2(din_04[2]),
  .ZN(_03954_)
);

NAND2_X1 _09460_ (
  .A1(_03952_),
  .A2(_03954_),
  .ZN(_03955_)
);

BUF_X2 _09461_ (
  .A(_03628_),
  .Z(_03956_)
);

NAND2_X1 _09462_ (
  .A1(_03955_),
  .A2(_03956_),
  .ZN(_03957_)
);

NAND2_X1 _09463_ (
  .A1(_03915_),
  .A2(\sresult[49][2] ),
  .ZN(_03958_)
);

NAND2_X1 _09464_ (
  .A1(_03957_),
  .A2(_03958_),
  .ZN(_00590_)
);

NAND2_X1 _09465_ (
  .A1(_03910_),
  .A2(\sresult[48][3] ),
  .ZN(_03959_)
);

NAND2_X1 _09466_ (
  .A1(_03953_),
  .A2(din_04[3]),
  .ZN(_03960_)
);

NAND2_X1 _09467_ (
  .A1(_03959_),
  .A2(_03960_),
  .ZN(_03961_)
);

NAND2_X1 _09468_ (
  .A1(_03961_),
  .A2(_03956_),
  .ZN(_03962_)
);

NAND2_X1 _09469_ (
  .A1(_03915_),
  .A2(\sresult[49][3] ),
  .ZN(_03963_)
);

NAND2_X1 _09470_ (
  .A1(_03962_),
  .A2(_03963_),
  .ZN(_00591_)
);

BUF_X4 _09471_ (
  .A(_03691_),
  .Z(_03964_)
);

NAND2_X1 _09472_ (
  .A1(_03964_),
  .A2(\sresult[48][4] ),
  .ZN(_03965_)
);

NAND2_X1 _09473_ (
  .A1(_03953_),
  .A2(din_04[4]),
  .ZN(_03966_)
);

NAND2_X1 _09474_ (
  .A1(_03965_),
  .A2(_03966_),
  .ZN(_03967_)
);

NAND2_X1 _09475_ (
  .A1(_03967_),
  .A2(_03956_),
  .ZN(_03968_)
);

BUF_X1 _09476_ (
  .A(_03752_),
  .Z(_03969_)
);

NAND2_X1 _09477_ (
  .A1(_03969_),
  .A2(\sresult[49][4] ),
  .ZN(_03970_)
);

NAND2_X1 _09478_ (
  .A1(_03968_),
  .A2(_03970_),
  .ZN(_00592_)
);

NAND2_X1 _09479_ (
  .A1(_03964_),
  .A2(\sresult[48][5] ),
  .ZN(_03971_)
);

NAND2_X1 _09480_ (
  .A1(_03953_),
  .A2(din_04[5]),
  .ZN(_03972_)
);

NAND2_X1 _09481_ (
  .A1(_03971_),
  .A2(_03972_),
  .ZN(_03973_)
);

NAND2_X1 _09482_ (
  .A1(_03973_),
  .A2(_03956_),
  .ZN(_03974_)
);

NAND2_X1 _09483_ (
  .A1(_03969_),
  .A2(\sresult[49][5] ),
  .ZN(_03975_)
);

NAND2_X1 _09484_ (
  .A1(_03974_),
  .A2(_03975_),
  .ZN(_00593_)
);

NAND2_X1 _09485_ (
  .A1(_03964_),
  .A2(\sresult[48][6] ),
  .ZN(_03976_)
);

NAND2_X1 _09486_ (
  .A1(_03953_),
  .A2(din_04[6]),
  .ZN(_03977_)
);

NAND2_X1 _09487_ (
  .A1(_03976_),
  .A2(_03977_),
  .ZN(_03978_)
);

NAND2_X1 _09488_ (
  .A1(_03978_),
  .A2(_03956_),
  .ZN(_03979_)
);

NAND2_X1 _09489_ (
  .A1(_03969_),
  .A2(\sresult[49][6] ),
  .ZN(_03980_)
);

NAND2_X1 _09490_ (
  .A1(_03979_),
  .A2(_03980_),
  .ZN(_00594_)
);

NAND2_X1 _09491_ (
  .A1(_03964_),
  .A2(\sresult[48][7] ),
  .ZN(_03981_)
);

NAND2_X1 _09492_ (
  .A1(_03953_),
  .A2(din_04[7]),
  .ZN(_03982_)
);

NAND2_X1 _09493_ (
  .A1(_03981_),
  .A2(_03982_),
  .ZN(_03983_)
);

NAND2_X1 _09494_ (
  .A1(_03983_),
  .A2(_03956_),
  .ZN(_03984_)
);

NAND2_X1 _09495_ (
  .A1(_03969_),
  .A2(\sresult[49][7] ),
  .ZN(_03985_)
);

NAND2_X1 _09496_ (
  .A1(_03984_),
  .A2(_03985_),
  .ZN(_00595_)
);

NAND2_X1 _09497_ (
  .A1(_03964_),
  .A2(\sresult[48][8] ),
  .ZN(_03986_)
);

NAND2_X1 _09498_ (
  .A1(_03953_),
  .A2(din_04[8]),
  .ZN(_03987_)
);

NAND2_X1 _09499_ (
  .A1(_03986_),
  .A2(_03987_),
  .ZN(_03988_)
);

NAND2_X1 _09500_ (
  .A1(_03988_),
  .A2(_03956_),
  .ZN(_03989_)
);

NAND2_X1 _09501_ (
  .A1(_03969_),
  .A2(\sresult[49][8] ),
  .ZN(_03990_)
);

NAND2_X1 _09502_ (
  .A1(_03989_),
  .A2(_03990_),
  .ZN(_00596_)
);

NAND2_X1 _09503_ (
  .A1(_03964_),
  .A2(\sresult[48][9] ),
  .ZN(_03991_)
);

NAND2_X1 _09504_ (
  .A1(_03953_),
  .A2(din_04[9]),
  .ZN(_03992_)
);

NAND2_X1 _09505_ (
  .A1(_03991_),
  .A2(_03992_),
  .ZN(_03993_)
);

NAND2_X1 _09506_ (
  .A1(_03993_),
  .A2(_03956_),
  .ZN(_03994_)
);

NAND2_X1 _09507_ (
  .A1(_03969_),
  .A2(\sresult[49][9] ),
  .ZN(_03995_)
);

NAND2_X1 _09508_ (
  .A1(_03994_),
  .A2(_03995_),
  .ZN(_00597_)
);

NAND2_X1 _09509_ (
  .A1(_03964_),
  .A2(\sresult[48][10] ),
  .ZN(_03996_)
);

NAND2_X1 _09510_ (
  .A1(_03953_),
  .A2(din_04[10]),
  .ZN(_03997_)
);

NAND2_X1 _09511_ (
  .A1(_03996_),
  .A2(_03997_),
  .ZN(_03998_)
);

NAND2_X1 _09512_ (
  .A1(_03998_),
  .A2(_03956_),
  .ZN(_03999_)
);

NAND2_X1 _09513_ (
  .A1(_03969_),
  .A2(\sresult[49][10] ),
  .ZN(_04000_)
);

NAND2_X1 _09514_ (
  .A1(_03999_),
  .A2(_04000_),
  .ZN(_00598_)
);

NAND2_X1 _09515_ (
  .A1(_03964_),
  .A2(\sresult[48][11] ),
  .ZN(_04001_)
);

NAND2_X1 _09516_ (
  .A1(_03953_),
  .A2(din_04[11]),
  .ZN(_04002_)
);

NAND2_X1 _09517_ (
  .A1(_04001_),
  .A2(_04002_),
  .ZN(_04003_)
);

NAND2_X1 _09518_ (
  .A1(_04003_),
  .A2(_03956_),
  .ZN(_04004_)
);

NAND2_X1 _09519_ (
  .A1(_03969_),
  .A2(\sresult[49][11] ),
  .ZN(_04005_)
);

NAND2_X1 _09520_ (
  .A1(_04004_),
  .A2(_04005_),
  .ZN(_00599_)
);

NAND2_X1 _09521_ (
  .A1(_03964_),
  .A2(\sresult[49][0] ),
  .ZN(_04006_)
);

BUF_X4 _09522_ (
  .A(_03735_),
  .Z(_04007_)
);

NAND2_X1 _09523_ (
  .A1(_04007_),
  .A2(din_13[0]),
  .ZN(_04008_)
);

NAND2_X1 _09524_ (
  .A1(_04006_),
  .A2(_04008_),
  .ZN(_04009_)
);

BUF_X2 _09525_ (
  .A(_03628_),
  .Z(_04010_)
);

NAND2_X1 _09526_ (
  .A1(_04009_),
  .A2(_04010_),
  .ZN(_04011_)
);

NAND2_X1 _09527_ (
  .A1(_03969_),
  .A2(\sresult[50][0] ),
  .ZN(_04012_)
);

NAND2_X1 _09528_ (
  .A1(_04011_),
  .A2(_04012_),
  .ZN(_00600_)
);

NAND2_X1 _09529_ (
  .A1(_03964_),
  .A2(\sresult[49][1] ),
  .ZN(_04013_)
);

NAND2_X1 _09530_ (
  .A1(_04007_),
  .A2(din_13[1]),
  .ZN(_04014_)
);

NAND2_X1 _09531_ (
  .A1(_04013_),
  .A2(_04014_),
  .ZN(_04015_)
);

NAND2_X1 _09532_ (
  .A1(_04015_),
  .A2(_04010_),
  .ZN(_04016_)
);

NAND2_X1 _09533_ (
  .A1(_03969_),
  .A2(\sresult[50][1] ),
  .ZN(_04017_)
);

NAND2_X1 _09534_ (
  .A1(_04016_),
  .A2(_04017_),
  .ZN(_00601_)
);

BUF_X4 _09535_ (
  .A(_03691_),
  .Z(_04018_)
);

NAND2_X1 _09536_ (
  .A1(_04018_),
  .A2(\sresult[49][2] ),
  .ZN(_04019_)
);

NAND2_X1 _09537_ (
  .A1(_04007_),
  .A2(din_13[2]),
  .ZN(_04020_)
);

NAND2_X1 _09538_ (
  .A1(_04019_),
  .A2(_04020_),
  .ZN(_04021_)
);

NAND2_X1 _09539_ (
  .A1(_04021_),
  .A2(_04010_),
  .ZN(_04022_)
);

BUF_X1 _09540_ (
  .A(_03752_),
  .Z(_04023_)
);

NAND2_X1 _09541_ (
  .A1(_04023_),
  .A2(\sresult[50][2] ),
  .ZN(_04024_)
);

NAND2_X1 _09542_ (
  .A1(_04022_),
  .A2(_04024_),
  .ZN(_00602_)
);

NAND2_X1 _09543_ (
  .A1(_04018_),
  .A2(\sresult[49][3] ),
  .ZN(_04025_)
);

NAND2_X1 _09544_ (
  .A1(_04007_),
  .A2(din_13[3]),
  .ZN(_04026_)
);

NAND2_X1 _09545_ (
  .A1(_04025_),
  .A2(_04026_),
  .ZN(_04027_)
);

NAND2_X1 _09546_ (
  .A1(_04027_),
  .A2(_04010_),
  .ZN(_04028_)
);

NAND2_X1 _09547_ (
  .A1(_04023_),
  .A2(\sresult[50][3] ),
  .ZN(_04029_)
);

NAND2_X1 _09548_ (
  .A1(_04028_),
  .A2(_04029_),
  .ZN(_00603_)
);

NAND2_X1 _09549_ (
  .A1(_04018_),
  .A2(\sresult[49][4] ),
  .ZN(_04030_)
);

NAND2_X1 _09550_ (
  .A1(_04007_),
  .A2(din_13[4]),
  .ZN(_04031_)
);

NAND2_X1 _09551_ (
  .A1(_04030_),
  .A2(_04031_),
  .ZN(_04032_)
);

NAND2_X1 _09552_ (
  .A1(_04032_),
  .A2(_04010_),
  .ZN(_04033_)
);

NAND2_X1 _09553_ (
  .A1(_04023_),
  .A2(\sresult[50][4] ),
  .ZN(_04034_)
);

NAND2_X1 _09554_ (
  .A1(_04033_),
  .A2(_04034_),
  .ZN(_00604_)
);

NAND2_X1 _09555_ (
  .A1(_04018_),
  .A2(\sresult[49][5] ),
  .ZN(_04035_)
);

NAND2_X1 _09556_ (
  .A1(_04007_),
  .A2(din_13[5]),
  .ZN(_04036_)
);

NAND2_X1 _09557_ (
  .A1(_04035_),
  .A2(_04036_),
  .ZN(_04037_)
);

NAND2_X1 _09558_ (
  .A1(_04037_),
  .A2(_04010_),
  .ZN(_04038_)
);

NAND2_X1 _09559_ (
  .A1(_04023_),
  .A2(\sresult[50][5] ),
  .ZN(_04039_)
);

NAND2_X1 _09560_ (
  .A1(_04038_),
  .A2(_04039_),
  .ZN(_00605_)
);

NAND2_X1 _09561_ (
  .A1(_04018_),
  .A2(\sresult[49][6] ),
  .ZN(_04040_)
);

NAND2_X1 _09562_ (
  .A1(_04007_),
  .A2(din_13[6]),
  .ZN(_04041_)
);

NAND2_X1 _09563_ (
  .A1(_04040_),
  .A2(_04041_),
  .ZN(_04042_)
);

NAND2_X1 _09564_ (
  .A1(_04042_),
  .A2(_04010_),
  .ZN(_04043_)
);

NAND2_X1 _09565_ (
  .A1(_04023_),
  .A2(\sresult[50][6] ),
  .ZN(_04044_)
);

NAND2_X1 _09566_ (
  .A1(_04043_),
  .A2(_04044_),
  .ZN(_00606_)
);

NAND2_X1 _09567_ (
  .A1(_04018_),
  .A2(\sresult[49][7] ),
  .ZN(_04045_)
);

NAND2_X1 _09568_ (
  .A1(_04007_),
  .A2(din_13[7]),
  .ZN(_04046_)
);

NAND2_X1 _09569_ (
  .A1(_04045_),
  .A2(_04046_),
  .ZN(_04047_)
);

NAND2_X1 _09570_ (
  .A1(_04047_),
  .A2(_04010_),
  .ZN(_04048_)
);

NAND2_X1 _09571_ (
  .A1(_04023_),
  .A2(\sresult[50][7] ),
  .ZN(_04049_)
);

NAND2_X1 _09572_ (
  .A1(_04048_),
  .A2(_04049_),
  .ZN(_00607_)
);

NAND2_X1 _09573_ (
  .A1(_04018_),
  .A2(\sresult[49][8] ),
  .ZN(_04050_)
);

NAND2_X1 _09574_ (
  .A1(_04007_),
  .A2(din_13[8]),
  .ZN(_04051_)
);

NAND2_X1 _09575_ (
  .A1(_04050_),
  .A2(_04051_),
  .ZN(_04052_)
);

NAND2_X1 _09576_ (
  .A1(_04052_),
  .A2(_04010_),
  .ZN(_04053_)
);

NAND2_X1 _09577_ (
  .A1(_04023_),
  .A2(\sresult[50][8] ),
  .ZN(_04054_)
);

NAND2_X1 _09578_ (
  .A1(_04053_),
  .A2(_04054_),
  .ZN(_00608_)
);

NAND2_X1 _09579_ (
  .A1(_04018_),
  .A2(\sresult[49][9] ),
  .ZN(_04055_)
);

NAND2_X1 _09580_ (
  .A1(_04007_),
  .A2(din_13[9]),
  .ZN(_04056_)
);

NAND2_X1 _09581_ (
  .A1(_04055_),
  .A2(_04056_),
  .ZN(_04057_)
);

NAND2_X1 _09582_ (
  .A1(_04057_),
  .A2(_04010_),
  .ZN(_04058_)
);

NAND2_X1 _09583_ (
  .A1(_04023_),
  .A2(\sresult[50][9] ),
  .ZN(_04059_)
);

NAND2_X1 _09584_ (
  .A1(_04058_),
  .A2(_04059_),
  .ZN(_00609_)
);

NAND2_X1 _09585_ (
  .A1(_04018_),
  .A2(\sresult[49][10] ),
  .ZN(_04060_)
);

BUF_X4 _09586_ (
  .A(_03735_),
  .Z(_04061_)
);

NAND2_X1 _09587_ (
  .A1(_04061_),
  .A2(din_13[10]),
  .ZN(_04062_)
);

NAND2_X1 _09588_ (
  .A1(_04060_),
  .A2(_04062_),
  .ZN(_04063_)
);

BUF_X2 _09589_ (
  .A(_03628_),
  .Z(_04064_)
);

NAND2_X1 _09590_ (
  .A1(_04063_),
  .A2(_04064_),
  .ZN(_04065_)
);

NAND2_X1 _09591_ (
  .A1(_04023_),
  .A2(\sresult[50][10] ),
  .ZN(_04066_)
);

NAND2_X1 _09592_ (
  .A1(_04065_),
  .A2(_04066_),
  .ZN(_00610_)
);

NAND2_X1 _09593_ (
  .A1(_04018_),
  .A2(\sresult[49][11] ),
  .ZN(_04067_)
);

NAND2_X1 _09594_ (
  .A1(_04061_),
  .A2(din_13[11]),
  .ZN(_04068_)
);

NAND2_X1 _09595_ (
  .A1(_04067_),
  .A2(_04068_),
  .ZN(_04069_)
);

NAND2_X1 _09596_ (
  .A1(_04069_),
  .A2(_04064_),
  .ZN(_04070_)
);

NAND2_X1 _09597_ (
  .A1(_04023_),
  .A2(\sresult[50][11] ),
  .ZN(_04071_)
);

NAND2_X1 _09598_ (
  .A1(_04070_),
  .A2(_04071_),
  .ZN(_00611_)
);

BUF_X4 _09599_ (
  .A(_03691_),
  .Z(_04072_)
);

NAND2_X1 _09600_ (
  .A1(_04072_),
  .A2(\sresult[50][0] ),
  .ZN(_04073_)
);

NAND2_X1 _09601_ (
  .A1(_04061_),
  .A2(din_22[0]),
  .ZN(_04074_)
);

NAND2_X1 _09602_ (
  .A1(_04073_),
  .A2(_04074_),
  .ZN(_04075_)
);

NAND2_X1 _09603_ (
  .A1(_04075_),
  .A2(_04064_),
  .ZN(_04076_)
);

BUF_X1 _09604_ (
  .A(_03752_),
  .Z(_04077_)
);

NAND2_X1 _09605_ (
  .A1(_04077_),
  .A2(\sresult[51][0] ),
  .ZN(_04078_)
);

NAND2_X1 _09606_ (
  .A1(_04076_),
  .A2(_04078_),
  .ZN(_00612_)
);

NAND2_X1 _09607_ (
  .A1(_04072_),
  .A2(\sresult[50][1] ),
  .ZN(_04079_)
);

NAND2_X1 _09608_ (
  .A1(_04061_),
  .A2(din_22[1]),
  .ZN(_04080_)
);

NAND2_X1 _09609_ (
  .A1(_04079_),
  .A2(_04080_),
  .ZN(_04081_)
);

NAND2_X1 _09610_ (
  .A1(_04081_),
  .A2(_04064_),
  .ZN(_04082_)
);

NAND2_X1 _09611_ (
  .A1(_04077_),
  .A2(\sresult[51][1] ),
  .ZN(_04083_)
);

NAND2_X1 _09612_ (
  .A1(_04082_),
  .A2(_04083_),
  .ZN(_00613_)
);

NAND2_X1 _09613_ (
  .A1(_04072_),
  .A2(\sresult[50][2] ),
  .ZN(_04084_)
);

NAND2_X1 _09614_ (
  .A1(_04061_),
  .A2(din_22[2]),
  .ZN(_04085_)
);

NAND2_X1 _09615_ (
  .A1(_04084_),
  .A2(_04085_),
  .ZN(_04086_)
);

NAND2_X1 _09616_ (
  .A1(_04086_),
  .A2(_04064_),
  .ZN(_04087_)
);

NAND2_X1 _09617_ (
  .A1(_04077_),
  .A2(\sresult[51][2] ),
  .ZN(_04088_)
);

NAND2_X1 _09618_ (
  .A1(_04087_),
  .A2(_04088_),
  .ZN(_00614_)
);

NAND2_X1 _09619_ (
  .A1(_04072_),
  .A2(\sresult[50][3] ),
  .ZN(_04089_)
);

NAND2_X1 _09620_ (
  .A1(_04061_),
  .A2(din_22[3]),
  .ZN(_04090_)
);

NAND2_X1 _09621_ (
  .A1(_04089_),
  .A2(_04090_),
  .ZN(_04091_)
);

NAND2_X1 _09622_ (
  .A1(_04091_),
  .A2(_04064_),
  .ZN(_04092_)
);

NAND2_X1 _09623_ (
  .A1(_04077_),
  .A2(\sresult[51][3] ),
  .ZN(_04093_)
);

NAND2_X1 _09624_ (
  .A1(_04092_),
  .A2(_04093_),
  .ZN(_00615_)
);

NAND2_X1 _09625_ (
  .A1(_04072_),
  .A2(\sresult[50][4] ),
  .ZN(_04094_)
);

NAND2_X1 _09626_ (
  .A1(_04061_),
  .A2(din_22[4]),
  .ZN(_04095_)
);

NAND2_X1 _09627_ (
  .A1(_04094_),
  .A2(_04095_),
  .ZN(_04096_)
);

NAND2_X1 _09628_ (
  .A1(_04096_),
  .A2(_04064_),
  .ZN(_04097_)
);

NAND2_X1 _09629_ (
  .A1(_04077_),
  .A2(\sresult[51][4] ),
  .ZN(_04098_)
);

NAND2_X1 _09630_ (
  .A1(_04097_),
  .A2(_04098_),
  .ZN(_00616_)
);

NAND2_X1 _09631_ (
  .A1(_04072_),
  .A2(\sresult[50][5] ),
  .ZN(_04099_)
);

NAND2_X1 _09632_ (
  .A1(_04061_),
  .A2(din_22[5]),
  .ZN(_04100_)
);

NAND2_X1 _09633_ (
  .A1(_04099_),
  .A2(_04100_),
  .ZN(_04101_)
);

NAND2_X1 _09634_ (
  .A1(_04101_),
  .A2(_04064_),
  .ZN(_04102_)
);

NAND2_X1 _09635_ (
  .A1(_04077_),
  .A2(\sresult[51][5] ),
  .ZN(_04103_)
);

NAND2_X1 _09636_ (
  .A1(_04102_),
  .A2(_04103_),
  .ZN(_00617_)
);

NAND2_X1 _09637_ (
  .A1(_04072_),
  .A2(\sresult[50][6] ),
  .ZN(_04104_)
);

NAND2_X1 _09638_ (
  .A1(_04061_),
  .A2(din_22[6]),
  .ZN(_04105_)
);

NAND2_X1 _09639_ (
  .A1(_04104_),
  .A2(_04105_),
  .ZN(_04106_)
);

NAND2_X1 _09640_ (
  .A1(_04106_),
  .A2(_04064_),
  .ZN(_04107_)
);

NAND2_X1 _09641_ (
  .A1(_04077_),
  .A2(\sresult[51][6] ),
  .ZN(_04108_)
);

NAND2_X1 _09642_ (
  .A1(_04107_),
  .A2(_04108_),
  .ZN(_00618_)
);

NAND2_X1 _09643_ (
  .A1(_04072_),
  .A2(\sresult[50][7] ),
  .ZN(_04109_)
);

NAND2_X1 _09644_ (
  .A1(_04061_),
  .A2(din_22[7]),
  .ZN(_04110_)
);

NAND2_X1 _09645_ (
  .A1(_04109_),
  .A2(_04110_),
  .ZN(_04111_)
);

NAND2_X1 _09646_ (
  .A1(_04111_),
  .A2(_04064_),
  .ZN(_04112_)
);

NAND2_X1 _09647_ (
  .A1(_04077_),
  .A2(\sresult[51][7] ),
  .ZN(_04113_)
);

NAND2_X1 _09648_ (
  .A1(_04112_),
  .A2(_04113_),
  .ZN(_00619_)
);

NAND2_X1 _09649_ (
  .A1(_04072_),
  .A2(\sresult[50][8] ),
  .ZN(_04114_)
);

BUF_X4 _09650_ (
  .A(_03735_),
  .Z(_04115_)
);

NAND2_X1 _09651_ (
  .A1(_04115_),
  .A2(din_22[8]),
  .ZN(_04116_)
);

NAND2_X1 _09652_ (
  .A1(_04114_),
  .A2(_04116_),
  .ZN(_04117_)
);

BUF_X2 _09653_ (
  .A(_03628_),
  .Z(_04118_)
);

NAND2_X1 _09654_ (
  .A1(_04117_),
  .A2(_04118_),
  .ZN(_04119_)
);

NAND2_X1 _09655_ (
  .A1(_04077_),
  .A2(\sresult[51][8] ),
  .ZN(_04120_)
);

NAND2_X1 _09656_ (
  .A1(_04119_),
  .A2(_04120_),
  .ZN(_00620_)
);

NAND2_X1 _09657_ (
  .A1(_04072_),
  .A2(\sresult[50][9] ),
  .ZN(_04121_)
);

NAND2_X1 _09658_ (
  .A1(_04115_),
  .A2(din_22[9]),
  .ZN(_04122_)
);

NAND2_X1 _09659_ (
  .A1(_04121_),
  .A2(_04122_),
  .ZN(_04123_)
);

NAND2_X1 _09660_ (
  .A1(_04123_),
  .A2(_04118_),
  .ZN(_04124_)
);

NAND2_X1 _09661_ (
  .A1(_04077_),
  .A2(\sresult[51][9] ),
  .ZN(_04125_)
);

NAND2_X1 _09662_ (
  .A1(_04124_),
  .A2(_04125_),
  .ZN(_00621_)
);

BUF_X4 _09663_ (
  .A(_03691_),
  .Z(_04126_)
);

NAND2_X1 _09664_ (
  .A1(_04126_),
  .A2(\sresult[50][10] ),
  .ZN(_04127_)
);

NAND2_X1 _09665_ (
  .A1(_04115_),
  .A2(din_22[10]),
  .ZN(_04128_)
);

NAND2_X1 _09666_ (
  .A1(_04127_),
  .A2(_04128_),
  .ZN(_04129_)
);

NAND2_X1 _09667_ (
  .A1(_04129_),
  .A2(_04118_),
  .ZN(_04130_)
);

BUF_X1 _09668_ (
  .A(_03752_),
  .Z(_04131_)
);

NAND2_X1 _09669_ (
  .A1(_04131_),
  .A2(\sresult[51][10] ),
  .ZN(_04132_)
);

NAND2_X1 _09670_ (
  .A1(_04130_),
  .A2(_04132_),
  .ZN(_00622_)
);

NAND2_X1 _09671_ (
  .A1(_04126_),
  .A2(\sresult[50][11] ),
  .ZN(_04133_)
);

NAND2_X1 _09672_ (
  .A1(_04115_),
  .A2(din_22[11]),
  .ZN(_04134_)
);

NAND2_X1 _09673_ (
  .A1(_04133_),
  .A2(_04134_),
  .ZN(_04135_)
);

NAND2_X1 _09674_ (
  .A1(_04135_),
  .A2(_04118_),
  .ZN(_04136_)
);

NAND2_X1 _09675_ (
  .A1(_04131_),
  .A2(\sresult[51][11] ),
  .ZN(_04137_)
);

NAND2_X1 _09676_ (
  .A1(_04136_),
  .A2(_04137_),
  .ZN(_00623_)
);

NAND2_X1 _09677_ (
  .A1(_04126_),
  .A2(\sresult[51][0] ),
  .ZN(_04138_)
);

NAND2_X1 _09678_ (
  .A1(_04115_),
  .A2(din_31[0]),
  .ZN(_04139_)
);

NAND2_X1 _09679_ (
  .A1(_04138_),
  .A2(_04139_),
  .ZN(_04140_)
);

NAND2_X1 _09680_ (
  .A1(_04140_),
  .A2(_04118_),
  .ZN(_04141_)
);

NAND2_X1 _09681_ (
  .A1(_04131_),
  .A2(\sresult[52][0] ),
  .ZN(_04142_)
);

NAND2_X1 _09682_ (
  .A1(_04141_),
  .A2(_04142_),
  .ZN(_00624_)
);

NAND2_X1 _09683_ (
  .A1(_04126_),
  .A2(\sresult[51][1] ),
  .ZN(_04143_)
);

NAND2_X1 _09684_ (
  .A1(_04115_),
  .A2(din_31[1]),
  .ZN(_04144_)
);

NAND2_X1 _09685_ (
  .A1(_04143_),
  .A2(_04144_),
  .ZN(_04145_)
);

NAND2_X1 _09686_ (
  .A1(_04145_),
  .A2(_04118_),
  .ZN(_04146_)
);

NAND2_X1 _09687_ (
  .A1(_04131_),
  .A2(\sresult[52][1] ),
  .ZN(_04147_)
);

NAND2_X1 _09688_ (
  .A1(_04146_),
  .A2(_04147_),
  .ZN(_00625_)
);

NAND2_X1 _09689_ (
  .A1(_04126_),
  .A2(\sresult[51][2] ),
  .ZN(_04148_)
);

NAND2_X1 _09690_ (
  .A1(_04115_),
  .A2(din_31[2]),
  .ZN(_04149_)
);

NAND2_X1 _09691_ (
  .A1(_04148_),
  .A2(_04149_),
  .ZN(_04150_)
);

NAND2_X1 _09692_ (
  .A1(_04150_),
  .A2(_04118_),
  .ZN(_04151_)
);

NAND2_X1 _09693_ (
  .A1(_04131_),
  .A2(\sresult[52][2] ),
  .ZN(_04152_)
);

NAND2_X1 _09694_ (
  .A1(_04151_),
  .A2(_04152_),
  .ZN(_00626_)
);

NAND2_X1 _09695_ (
  .A1(_04126_),
  .A2(\sresult[51][3] ),
  .ZN(_04153_)
);

NAND2_X1 _09696_ (
  .A1(_04115_),
  .A2(din_31[3]),
  .ZN(_04154_)
);

NAND2_X1 _09697_ (
  .A1(_04153_),
  .A2(_04154_),
  .ZN(_04155_)
);

NAND2_X1 _09698_ (
  .A1(_04155_),
  .A2(_04118_),
  .ZN(_04156_)
);

NAND2_X1 _09699_ (
  .A1(_04131_),
  .A2(\sresult[52][3] ),
  .ZN(_04157_)
);

NAND2_X1 _09700_ (
  .A1(_04156_),
  .A2(_04157_),
  .ZN(_00627_)
);

NAND2_X1 _09701_ (
  .A1(_04126_),
  .A2(\sresult[51][4] ),
  .ZN(_04158_)
);

NAND2_X1 _09702_ (
  .A1(_04115_),
  .A2(din_31[4]),
  .ZN(_04159_)
);

NAND2_X1 _09703_ (
  .A1(_04158_),
  .A2(_04159_),
  .ZN(_04160_)
);

NAND2_X1 _09704_ (
  .A1(_04160_),
  .A2(_04118_),
  .ZN(_04161_)
);

NAND2_X1 _09705_ (
  .A1(_04131_),
  .A2(\sresult[52][4] ),
  .ZN(_04162_)
);

NAND2_X1 _09706_ (
  .A1(_04161_),
  .A2(_04162_),
  .ZN(_00628_)
);

NAND2_X1 _09707_ (
  .A1(_04126_),
  .A2(\sresult[51][5] ),
  .ZN(_04163_)
);

NAND2_X1 _09708_ (
  .A1(_04115_),
  .A2(din_31[5]),
  .ZN(_04164_)
);

NAND2_X1 _09709_ (
  .A1(_04163_),
  .A2(_04164_),
  .ZN(_04165_)
);

NAND2_X1 _09710_ (
  .A1(_04165_),
  .A2(_04118_),
  .ZN(_04166_)
);

NAND2_X1 _09711_ (
  .A1(_04131_),
  .A2(\sresult[52][5] ),
  .ZN(_04167_)
);

NAND2_X1 _09712_ (
  .A1(_04166_),
  .A2(_04167_),
  .ZN(_00629_)
);

NAND2_X1 _09713_ (
  .A1(_04126_),
  .A2(\sresult[51][6] ),
  .ZN(_04168_)
);

BUF_X4 _09714_ (
  .A(_03735_),
  .Z(_04169_)
);

NAND2_X1 _09715_ (
  .A1(_04169_),
  .A2(din_31[6]),
  .ZN(_04170_)
);

NAND2_X1 _09716_ (
  .A1(_04168_),
  .A2(_04170_),
  .ZN(_04171_)
);

BUF_X4 _09717_ (
  .A(_00911_),
  .Z(_04172_)
);

BUF_X2 _09718_ (
  .A(_04172_),
  .Z(_04173_)
);

NAND2_X1 _09719_ (
  .A1(_04171_),
  .A2(_04173_),
  .ZN(_04174_)
);

NAND2_X1 _09720_ (
  .A1(_04131_),
  .A2(\sresult[52][6] ),
  .ZN(_04175_)
);

NAND2_X1 _09721_ (
  .A1(_04174_),
  .A2(_04175_),
  .ZN(_00630_)
);

NAND2_X1 _09722_ (
  .A1(_04126_),
  .A2(\sresult[51][7] ),
  .ZN(_04176_)
);

NAND2_X1 _09723_ (
  .A1(_04169_),
  .A2(din_31[7]),
  .ZN(_04177_)
);

NAND2_X1 _09724_ (
  .A1(_04176_),
  .A2(_04177_),
  .ZN(_04178_)
);

NAND2_X1 _09725_ (
  .A1(_04178_),
  .A2(_04173_),
  .ZN(_04179_)
);

NAND2_X1 _09726_ (
  .A1(_04131_),
  .A2(\sresult[52][7] ),
  .ZN(_04180_)
);

NAND2_X1 _09727_ (
  .A1(_04179_),
  .A2(_04180_),
  .ZN(_00631_)
);

BUF_X4 _09728_ (
  .A(_03691_),
  .Z(_04181_)
);

NAND2_X1 _09729_ (
  .A1(_04181_),
  .A2(\sresult[51][8] ),
  .ZN(_04182_)
);

NAND2_X1 _09730_ (
  .A1(_04169_),
  .A2(din_31[8]),
  .ZN(_04183_)
);

NAND2_X1 _09731_ (
  .A1(_04182_),
  .A2(_04183_),
  .ZN(_04184_)
);

NAND2_X1 _09732_ (
  .A1(_04184_),
  .A2(_04173_),
  .ZN(_04185_)
);

BUF_X1 _09733_ (
  .A(_03752_),
  .Z(_04186_)
);

NAND2_X1 _09734_ (
  .A1(_04186_),
  .A2(\sresult[52][8] ),
  .ZN(_04187_)
);

NAND2_X1 _09735_ (
  .A1(_04185_),
  .A2(_04187_),
  .ZN(_00632_)
);

NAND2_X1 _09736_ (
  .A1(_04181_),
  .A2(\sresult[51][9] ),
  .ZN(_04188_)
);

NAND2_X1 _09737_ (
  .A1(_04169_),
  .A2(din_31[9]),
  .ZN(_04189_)
);

NAND2_X1 _09738_ (
  .A1(_04188_),
  .A2(_04189_),
  .ZN(_04190_)
);

NAND2_X1 _09739_ (
  .A1(_04190_),
  .A2(_04173_),
  .ZN(_04191_)
);

NAND2_X1 _09740_ (
  .A1(_04186_),
  .A2(\sresult[52][9] ),
  .ZN(_04192_)
);

NAND2_X1 _09741_ (
  .A1(_04191_),
  .A2(_04192_),
  .ZN(_00633_)
);

NAND2_X1 _09742_ (
  .A1(_04181_),
  .A2(\sresult[51][10] ),
  .ZN(_04193_)
);

NAND2_X1 _09743_ (
  .A1(_04169_),
  .A2(din_31[10]),
  .ZN(_04194_)
);

NAND2_X1 _09744_ (
  .A1(_04193_),
  .A2(_04194_),
  .ZN(_04195_)
);

NAND2_X1 _09745_ (
  .A1(_04195_),
  .A2(_04173_),
  .ZN(_04196_)
);

NAND2_X1 _09746_ (
  .A1(_04186_),
  .A2(\sresult[52][10] ),
  .ZN(_04197_)
);

NAND2_X1 _09747_ (
  .A1(_04196_),
  .A2(_04197_),
  .ZN(_00634_)
);

NAND2_X1 _09748_ (
  .A1(_04181_),
  .A2(\sresult[51][11] ),
  .ZN(_04198_)
);

NAND2_X1 _09749_ (
  .A1(_04169_),
  .A2(din_31[11]),
  .ZN(_04199_)
);

NAND2_X1 _09750_ (
  .A1(_04198_),
  .A2(_04199_),
  .ZN(_04200_)
);

NAND2_X1 _09751_ (
  .A1(_04200_),
  .A2(_04173_),
  .ZN(_04201_)
);

NAND2_X1 _09752_ (
  .A1(_04186_),
  .A2(\sresult[52][11] ),
  .ZN(_04202_)
);

NAND2_X1 _09753_ (
  .A1(_04201_),
  .A2(_04202_),
  .ZN(_00635_)
);

NAND2_X1 _09754_ (
  .A1(_04181_),
  .A2(\sresult[52][0] ),
  .ZN(_04203_)
);

NAND2_X1 _09755_ (
  .A1(_04169_),
  .A2(din_40[0]),
  .ZN(_04204_)
);

NAND2_X1 _09756_ (
  .A1(_04203_),
  .A2(_04204_),
  .ZN(_04205_)
);

NAND2_X1 _09757_ (
  .A1(_04205_),
  .A2(_04173_),
  .ZN(_04206_)
);

NAND2_X1 _09758_ (
  .A1(_04186_),
  .A2(\sresult[53][0] ),
  .ZN(_04207_)
);

NAND2_X1 _09759_ (
  .A1(_04206_),
  .A2(_04207_),
  .ZN(_00636_)
);

NAND2_X1 _09760_ (
  .A1(_04181_),
  .A2(\sresult[52][1] ),
  .ZN(_04208_)
);

NAND2_X1 _09761_ (
  .A1(_04169_),
  .A2(din_40[1]),
  .ZN(_04209_)
);

NAND2_X1 _09762_ (
  .A1(_04208_),
  .A2(_04209_),
  .ZN(_04210_)
);

NAND2_X1 _09763_ (
  .A1(_04210_),
  .A2(_04173_),
  .ZN(_04211_)
);

NAND2_X1 _09764_ (
  .A1(_04186_),
  .A2(\sresult[53][1] ),
  .ZN(_04212_)
);

NAND2_X1 _09765_ (
  .A1(_04211_),
  .A2(_04212_),
  .ZN(_00637_)
);

NAND2_X1 _09766_ (
  .A1(_04181_),
  .A2(\sresult[52][2] ),
  .ZN(_04213_)
);

NAND2_X1 _09767_ (
  .A1(_04169_),
  .A2(din_40[2]),
  .ZN(_04214_)
);

NAND2_X1 _09768_ (
  .A1(_04213_),
  .A2(_04214_),
  .ZN(_04215_)
);

NAND2_X1 _09769_ (
  .A1(_04215_),
  .A2(_04173_),
  .ZN(_04216_)
);

NAND2_X1 _09770_ (
  .A1(_04186_),
  .A2(\sresult[53][2] ),
  .ZN(_04217_)
);

NAND2_X1 _09771_ (
  .A1(_04216_),
  .A2(_04217_),
  .ZN(_00638_)
);

NAND2_X1 _09772_ (
  .A1(_04181_),
  .A2(\sresult[52][3] ),
  .ZN(_04218_)
);

NAND2_X1 _09773_ (
  .A1(_04169_),
  .A2(din_40[3]),
  .ZN(_04219_)
);

NAND2_X1 _09774_ (
  .A1(_04218_),
  .A2(_04219_),
  .ZN(_04220_)
);

NAND2_X1 _09775_ (
  .A1(_04220_),
  .A2(_04173_),
  .ZN(_04221_)
);

NAND2_X1 _09776_ (
  .A1(_04186_),
  .A2(\sresult[53][3] ),
  .ZN(_04222_)
);

NAND2_X1 _09777_ (
  .A1(_04221_),
  .A2(_04222_),
  .ZN(_00639_)
);

NAND2_X1 _09778_ (
  .A1(_04181_),
  .A2(\sresult[52][4] ),
  .ZN(_04223_)
);

BUF_X4 _09779_ (
  .A(_03735_),
  .Z(_04224_)
);

NAND2_X1 _09780_ (
  .A1(_04224_),
  .A2(din_40[4]),
  .ZN(_04225_)
);

NAND2_X1 _09781_ (
  .A1(_04223_),
  .A2(_04225_),
  .ZN(_04226_)
);

BUF_X2 _09782_ (
  .A(_04172_),
  .Z(_04227_)
);

NAND2_X1 _09783_ (
  .A1(_04226_),
  .A2(_04227_),
  .ZN(_04228_)
);

NAND2_X1 _09784_ (
  .A1(_04186_),
  .A2(\sresult[53][4] ),
  .ZN(_04229_)
);

NAND2_X1 _09785_ (
  .A1(_04228_),
  .A2(_04229_),
  .ZN(_00640_)
);

NAND2_X1 _09786_ (
  .A1(_04181_),
  .A2(\sresult[52][5] ),
  .ZN(_04230_)
);

NAND2_X1 _09787_ (
  .A1(_04224_),
  .A2(din_40[5]),
  .ZN(_04231_)
);

NAND2_X1 _09788_ (
  .A1(_04230_),
  .A2(_04231_),
  .ZN(_04232_)
);

NAND2_X1 _09789_ (
  .A1(_04232_),
  .A2(_04227_),
  .ZN(_04233_)
);

NAND2_X1 _09790_ (
  .A1(_04186_),
  .A2(\sresult[53][5] ),
  .ZN(_04234_)
);

NAND2_X1 _09791_ (
  .A1(_04233_),
  .A2(_04234_),
  .ZN(_00641_)
);

BUF_X8 _09792_ (
  .A(_00799_),
  .Z(_04235_)
);

BUF_X4 _09793_ (
  .A(_04235_),
  .Z(_04236_)
);

NAND2_X1 _09794_ (
  .A1(_04236_),
  .A2(\sresult[52][6] ),
  .ZN(_04237_)
);

NAND2_X1 _09795_ (
  .A1(_04224_),
  .A2(din_40[6]),
  .ZN(_04238_)
);

NAND2_X1 _09796_ (
  .A1(_04237_),
  .A2(_04238_),
  .ZN(_04239_)
);

NAND2_X1 _09797_ (
  .A1(_04239_),
  .A2(_04227_),
  .ZN(_04240_)
);

BUF_X1 _09798_ (
  .A(_03752_),
  .Z(_04241_)
);

NAND2_X1 _09799_ (
  .A1(_04241_),
  .A2(\sresult[53][6] ),
  .ZN(_04242_)
);

NAND2_X1 _09800_ (
  .A1(_04240_),
  .A2(_04242_),
  .ZN(_00642_)
);

NAND2_X1 _09801_ (
  .A1(_04236_),
  .A2(\sresult[52][7] ),
  .ZN(_04243_)
);

NAND2_X1 _09802_ (
  .A1(_04224_),
  .A2(din_40[7]),
  .ZN(_04244_)
);

NAND2_X1 _09803_ (
  .A1(_04243_),
  .A2(_04244_),
  .ZN(_04245_)
);

NAND2_X1 _09804_ (
  .A1(_04245_),
  .A2(_04227_),
  .ZN(_04246_)
);

NAND2_X1 _09805_ (
  .A1(_04241_),
  .A2(\sresult[53][7] ),
  .ZN(_04247_)
);

NAND2_X1 _09806_ (
  .A1(_04246_),
  .A2(_04247_),
  .ZN(_00643_)
);

NAND2_X1 _09807_ (
  .A1(_04236_),
  .A2(\sresult[52][8] ),
  .ZN(_04248_)
);

NAND2_X1 _09808_ (
  .A1(_04224_),
  .A2(din_40[8]),
  .ZN(_04249_)
);

NAND2_X1 _09809_ (
  .A1(_04248_),
  .A2(_04249_),
  .ZN(_04250_)
);

NAND2_X1 _09810_ (
  .A1(_04250_),
  .A2(_04227_),
  .ZN(_04251_)
);

NAND2_X1 _09811_ (
  .A1(_04241_),
  .A2(\sresult[53][8] ),
  .ZN(_04252_)
);

NAND2_X1 _09812_ (
  .A1(_04251_),
  .A2(_04252_),
  .ZN(_00644_)
);

NAND2_X1 _09813_ (
  .A1(_04236_),
  .A2(\sresult[52][9] ),
  .ZN(_04253_)
);

NAND2_X1 _09814_ (
  .A1(_04224_),
  .A2(din_40[9]),
  .ZN(_04254_)
);

NAND2_X1 _09815_ (
  .A1(_04253_),
  .A2(_04254_),
  .ZN(_04255_)
);

NAND2_X1 _09816_ (
  .A1(_04255_),
  .A2(_04227_),
  .ZN(_04256_)
);

NAND2_X1 _09817_ (
  .A1(_04241_),
  .A2(\sresult[53][9] ),
  .ZN(_04257_)
);

NAND2_X1 _09818_ (
  .A1(_04256_),
  .A2(_04257_),
  .ZN(_00645_)
);

NAND2_X1 _09819_ (
  .A1(_04236_),
  .A2(\sresult[52][10] ),
  .ZN(_04258_)
);

NAND2_X1 _09820_ (
  .A1(_04224_),
  .A2(din_40[10]),
  .ZN(_04259_)
);

NAND2_X1 _09821_ (
  .A1(_04258_),
  .A2(_04259_),
  .ZN(_04260_)
);

NAND2_X1 _09822_ (
  .A1(_04260_),
  .A2(_04227_),
  .ZN(_04261_)
);

NAND2_X1 _09823_ (
  .A1(_04241_),
  .A2(\sresult[53][10] ),
  .ZN(_04262_)
);

NAND2_X1 _09824_ (
  .A1(_04261_),
  .A2(_04262_),
  .ZN(_00646_)
);

NAND2_X1 _09825_ (
  .A1(_04236_),
  .A2(\sresult[52][11] ),
  .ZN(_04263_)
);

NAND2_X1 _09826_ (
  .A1(_04224_),
  .A2(din_40[11]),
  .ZN(_04264_)
);

NAND2_X1 _09827_ (
  .A1(_04263_),
  .A2(_04264_),
  .ZN(_04265_)
);

NAND2_X1 _09828_ (
  .A1(_04265_),
  .A2(_04227_),
  .ZN(_04266_)
);

NAND2_X1 _09829_ (
  .A1(_04241_),
  .A2(\sresult[53][11] ),
  .ZN(_04267_)
);

NAND2_X1 _09830_ (
  .A1(_04266_),
  .A2(_04267_),
  .ZN(_00647_)
);

NAND2_X1 _09831_ (
  .A1(_04236_),
  .A2(\sresult[53][0] ),
  .ZN(_04268_)
);

NAND2_X1 _09832_ (
  .A1(_04224_),
  .A2(din_30[0]),
  .ZN(_04269_)
);

NAND2_X1 _09833_ (
  .A1(_04268_),
  .A2(_04269_),
  .ZN(_04270_)
);

NAND2_X1 _09834_ (
  .A1(_04270_),
  .A2(_04227_),
  .ZN(_04271_)
);

NAND2_X1 _09835_ (
  .A1(_04241_),
  .A2(\sresult[54][0] ),
  .ZN(_04272_)
);

NAND2_X1 _09836_ (
  .A1(_04271_),
  .A2(_04272_),
  .ZN(_00648_)
);

NAND2_X1 _09837_ (
  .A1(_04236_),
  .A2(\sresult[53][1] ),
  .ZN(_04273_)
);

NAND2_X1 _09838_ (
  .A1(_04224_),
  .A2(din_30[1]),
  .ZN(_04274_)
);

NAND2_X1 _09839_ (
  .A1(_04273_),
  .A2(_04274_),
  .ZN(_04275_)
);

NAND2_X1 _09840_ (
  .A1(_04275_),
  .A2(_04227_),
  .ZN(_04276_)
);

NAND2_X1 _09841_ (
  .A1(_04241_),
  .A2(\sresult[54][1] ),
  .ZN(_04277_)
);

NAND2_X1 _09842_ (
  .A1(_04276_),
  .A2(_04277_),
  .ZN(_00649_)
);

NAND2_X1 _09843_ (
  .A1(_04236_),
  .A2(\sresult[53][2] ),
  .ZN(_04278_)
);

BUF_X8 _09844_ (
  .A(_00770_),
  .Z(_04279_)
);

BUF_X4 _09845_ (
  .A(_04279_),
  .Z(_04280_)
);

NAND2_X1 _09846_ (
  .A1(_04280_),
  .A2(din_30[2]),
  .ZN(_04281_)
);

NAND2_X1 _09847_ (
  .A1(_04278_),
  .A2(_04281_),
  .ZN(_04282_)
);

BUF_X2 _09848_ (
  .A(_04172_),
  .Z(_04283_)
);

NAND2_X1 _09849_ (
  .A1(_04282_),
  .A2(_04283_),
  .ZN(_04284_)
);

NAND2_X1 _09850_ (
  .A1(_04241_),
  .A2(\sresult[54][2] ),
  .ZN(_04285_)
);

NAND2_X1 _09851_ (
  .A1(_04284_),
  .A2(_04285_),
  .ZN(_00650_)
);

NAND2_X1 _09852_ (
  .A1(_04236_),
  .A2(\sresult[53][3] ),
  .ZN(_04286_)
);

NAND2_X1 _09853_ (
  .A1(_04280_),
  .A2(din_30[3]),
  .ZN(_04287_)
);

NAND2_X1 _09854_ (
  .A1(_04286_),
  .A2(_04287_),
  .ZN(_04288_)
);

NAND2_X1 _09855_ (
  .A1(_04288_),
  .A2(_04283_),
  .ZN(_04289_)
);

NAND2_X1 _09856_ (
  .A1(_04241_),
  .A2(\sresult[54][3] ),
  .ZN(_04290_)
);

NAND2_X1 _09857_ (
  .A1(_04289_),
  .A2(_04290_),
  .ZN(_00651_)
);

BUF_X4 _09858_ (
  .A(_04235_),
  .Z(_04291_)
);

NAND2_X1 _09859_ (
  .A1(_04291_),
  .A2(\sresult[53][4] ),
  .ZN(_04292_)
);

NAND2_X1 _09860_ (
  .A1(_04280_),
  .A2(din_30[4]),
  .ZN(_04293_)
);

NAND2_X1 _09861_ (
  .A1(_04292_),
  .A2(_04293_),
  .ZN(_04294_)
);

NAND2_X1 _09862_ (
  .A1(_04294_),
  .A2(_04283_),
  .ZN(_04295_)
);

BUF_X4 _09863_ (
  .A(_00810_),
  .Z(_04296_)
);

CLKBUF_X2 _09864_ (
  .A(_04296_),
  .Z(_04297_)
);

NAND2_X1 _09865_ (
  .A1(_04297_),
  .A2(\sresult[54][4] ),
  .ZN(_04298_)
);

NAND2_X1 _09866_ (
  .A1(_04295_),
  .A2(_04298_),
  .ZN(_00652_)
);

NAND2_X1 _09867_ (
  .A1(_04291_),
  .A2(\sresult[53][5] ),
  .ZN(_04299_)
);

NAND2_X1 _09868_ (
  .A1(_04280_),
  .A2(din_30[5]),
  .ZN(_04300_)
);

NAND2_X1 _09869_ (
  .A1(_04299_),
  .A2(_04300_),
  .ZN(_04301_)
);

NAND2_X1 _09870_ (
  .A1(_04301_),
  .A2(_04283_),
  .ZN(_04302_)
);

NAND2_X1 _09871_ (
  .A1(_04297_),
  .A2(\sresult[54][5] ),
  .ZN(_04303_)
);

NAND2_X1 _09872_ (
  .A1(_04302_),
  .A2(_04303_),
  .ZN(_00653_)
);

NAND2_X1 _09873_ (
  .A1(_04291_),
  .A2(\sresult[53][6] ),
  .ZN(_04304_)
);

NAND2_X1 _09874_ (
  .A1(_04280_),
  .A2(din_30[6]),
  .ZN(_04305_)
);

NAND2_X1 _09875_ (
  .A1(_04304_),
  .A2(_04305_),
  .ZN(_04306_)
);

NAND2_X1 _09876_ (
  .A1(_04306_),
  .A2(_04283_),
  .ZN(_04307_)
);

NAND2_X1 _09877_ (
  .A1(_04297_),
  .A2(\sresult[54][6] ),
  .ZN(_04308_)
);

NAND2_X1 _09878_ (
  .A1(_04307_),
  .A2(_04308_),
  .ZN(_00654_)
);

NAND2_X1 _09879_ (
  .A1(_04291_),
  .A2(\sresult[53][7] ),
  .ZN(_04309_)
);

NAND2_X1 _09880_ (
  .A1(_04280_),
  .A2(din_30[7]),
  .ZN(_04310_)
);

NAND2_X1 _09881_ (
  .A1(_04309_),
  .A2(_04310_),
  .ZN(_04311_)
);

NAND2_X1 _09882_ (
  .A1(_04311_),
  .A2(_04283_),
  .ZN(_04312_)
);

NAND2_X1 _09883_ (
  .A1(_04297_),
  .A2(\sresult[54][7] ),
  .ZN(_04313_)
);

NAND2_X1 _09884_ (
  .A1(_04312_),
  .A2(_04313_),
  .ZN(_00655_)
);

NAND2_X1 _09885_ (
  .A1(_04291_),
  .A2(\sresult[53][8] ),
  .ZN(_04314_)
);

NAND2_X1 _09886_ (
  .A1(_04280_),
  .A2(din_30[8]),
  .ZN(_04315_)
);

NAND2_X1 _09887_ (
  .A1(_04314_),
  .A2(_04315_),
  .ZN(_04316_)
);

NAND2_X1 _09888_ (
  .A1(_04316_),
  .A2(_04283_),
  .ZN(_04317_)
);

NAND2_X1 _09889_ (
  .A1(_04297_),
  .A2(\sresult[54][8] ),
  .ZN(_04318_)
);

NAND2_X1 _09890_ (
  .A1(_04317_),
  .A2(_04318_),
  .ZN(_00656_)
);

NAND2_X1 _09891_ (
  .A1(_04291_),
  .A2(\sresult[53][9] ),
  .ZN(_04319_)
);

NAND2_X1 _09892_ (
  .A1(_04280_),
  .A2(din_30[9]),
  .ZN(_04320_)
);

NAND2_X1 _09893_ (
  .A1(_04319_),
  .A2(_04320_),
  .ZN(_04321_)
);

NAND2_X1 _09894_ (
  .A1(_04321_),
  .A2(_04283_),
  .ZN(_04322_)
);

NAND2_X1 _09895_ (
  .A1(_04297_),
  .A2(\sresult[54][9] ),
  .ZN(_04323_)
);

NAND2_X1 _09896_ (
  .A1(_04322_),
  .A2(_04323_),
  .ZN(_00657_)
);

NAND2_X1 _09897_ (
  .A1(_04291_),
  .A2(\sresult[53][10] ),
  .ZN(_04324_)
);

NAND2_X1 _09898_ (
  .A1(_04280_),
  .A2(din_30[10]),
  .ZN(_04325_)
);

NAND2_X1 _09899_ (
  .A1(_04324_),
  .A2(_04325_),
  .ZN(_04326_)
);

NAND2_X1 _09900_ (
  .A1(_04326_),
  .A2(_04283_),
  .ZN(_04327_)
);

NAND2_X1 _09901_ (
  .A1(_04297_),
  .A2(\sresult[54][10] ),
  .ZN(_04328_)
);

NAND2_X1 _09902_ (
  .A1(_04327_),
  .A2(_04328_),
  .ZN(_00658_)
);

NAND2_X1 _09903_ (
  .A1(_04291_),
  .A2(\sresult[53][11] ),
  .ZN(_04329_)
);

NAND2_X1 _09904_ (
  .A1(_04280_),
  .A2(din_30[11]),
  .ZN(_04330_)
);

NAND2_X1 _09905_ (
  .A1(_04329_),
  .A2(_04330_),
  .ZN(_04331_)
);

NAND2_X1 _09906_ (
  .A1(_04331_),
  .A2(_04283_),
  .ZN(_04332_)
);

NAND2_X1 _09907_ (
  .A1(_04297_),
  .A2(\sresult[54][11] ),
  .ZN(_04333_)
);

NAND2_X1 _09908_ (
  .A1(_04332_),
  .A2(_04333_),
  .ZN(_00659_)
);

NAND2_X1 _09909_ (
  .A1(_04291_),
  .A2(\sresult[54][0] ),
  .ZN(_04334_)
);

BUF_X4 _09910_ (
  .A(_04279_),
  .Z(_04335_)
);

NAND2_X1 _09911_ (
  .A1(_04335_),
  .A2(din_21[0]),
  .ZN(_04336_)
);

NAND2_X1 _09912_ (
  .A1(_04334_),
  .A2(_04336_),
  .ZN(_04337_)
);

BUF_X2 _09913_ (
  .A(_04172_),
  .Z(_04338_)
);

NAND2_X1 _09914_ (
  .A1(_04337_),
  .A2(_04338_),
  .ZN(_04339_)
);

NAND2_X1 _09915_ (
  .A1(_04297_),
  .A2(\sresult[55][0] ),
  .ZN(_04340_)
);

NAND2_X1 _09916_ (
  .A1(_04339_),
  .A2(_04340_),
  .ZN(_00660_)
);

NAND2_X1 _09917_ (
  .A1(_04291_),
  .A2(\sresult[54][1] ),
  .ZN(_04341_)
);

NAND2_X1 _09918_ (
  .A1(_04335_),
  .A2(din_21[1]),
  .ZN(_04342_)
);

NAND2_X1 _09919_ (
  .A1(_04341_),
  .A2(_04342_),
  .ZN(_04343_)
);

NAND2_X1 _09920_ (
  .A1(_04343_),
  .A2(_04338_),
  .ZN(_04344_)
);

NAND2_X1 _09921_ (
  .A1(_04297_),
  .A2(\sresult[55][1] ),
  .ZN(_04345_)
);

NAND2_X1 _09922_ (
  .A1(_04344_),
  .A2(_04345_),
  .ZN(_00661_)
);

BUF_X4 _09923_ (
  .A(_04235_),
  .Z(_04346_)
);

NAND2_X1 _09924_ (
  .A1(_04346_),
  .A2(\sresult[54][2] ),
  .ZN(_04347_)
);

NAND2_X1 _09925_ (
  .A1(_04335_),
  .A2(din_21[2]),
  .ZN(_04348_)
);

NAND2_X1 _09926_ (
  .A1(_04347_),
  .A2(_04348_),
  .ZN(_04349_)
);

NAND2_X1 _09927_ (
  .A1(_04349_),
  .A2(_04338_),
  .ZN(_04350_)
);

CLKBUF_X2 _09928_ (
  .A(_04296_),
  .Z(_04351_)
);

NAND2_X1 _09929_ (
  .A1(_04351_),
  .A2(\sresult[55][2] ),
  .ZN(_04352_)
);

NAND2_X1 _09930_ (
  .A1(_04350_),
  .A2(_04352_),
  .ZN(_00662_)
);

NAND2_X1 _09931_ (
  .A1(_04346_),
  .A2(\sresult[54][3] ),
  .ZN(_04353_)
);

NAND2_X1 _09932_ (
  .A1(_04335_),
  .A2(din_21[3]),
  .ZN(_04354_)
);

NAND2_X1 _09933_ (
  .A1(_04353_),
  .A2(_04354_),
  .ZN(_04355_)
);

NAND2_X1 _09934_ (
  .A1(_04355_),
  .A2(_04338_),
  .ZN(_04356_)
);

NAND2_X1 _09935_ (
  .A1(_04351_),
  .A2(\sresult[55][3] ),
  .ZN(_04357_)
);

NAND2_X1 _09936_ (
  .A1(_04356_),
  .A2(_04357_),
  .ZN(_00663_)
);

NAND2_X1 _09937_ (
  .A1(_04346_),
  .A2(\sresult[54][4] ),
  .ZN(_04358_)
);

NAND2_X1 _09938_ (
  .A1(_04335_),
  .A2(din_21[4]),
  .ZN(_04359_)
);

NAND2_X1 _09939_ (
  .A1(_04358_),
  .A2(_04359_),
  .ZN(_04360_)
);

NAND2_X1 _09940_ (
  .A1(_04360_),
  .A2(_04338_),
  .ZN(_04361_)
);

NAND2_X1 _09941_ (
  .A1(_04351_),
  .A2(\sresult[55][4] ),
  .ZN(_04362_)
);

NAND2_X1 _09942_ (
  .A1(_04361_),
  .A2(_04362_),
  .ZN(_00664_)
);

NAND2_X1 _09943_ (
  .A1(_04346_),
  .A2(\sresult[54][5] ),
  .ZN(_04363_)
);

NAND2_X1 _09944_ (
  .A1(_04335_),
  .A2(din_21[5]),
  .ZN(_04364_)
);

NAND2_X1 _09945_ (
  .A1(_04363_),
  .A2(_04364_),
  .ZN(_04365_)
);

NAND2_X1 _09946_ (
  .A1(_04365_),
  .A2(_04338_),
  .ZN(_04366_)
);

NAND2_X1 _09947_ (
  .A1(_04351_),
  .A2(\sresult[55][5] ),
  .ZN(_04367_)
);

NAND2_X1 _09948_ (
  .A1(_04366_),
  .A2(_04367_),
  .ZN(_00665_)
);

NAND2_X1 _09949_ (
  .A1(_04346_),
  .A2(\sresult[54][6] ),
  .ZN(_04368_)
);

NAND2_X1 _09950_ (
  .A1(_04335_),
  .A2(din_21[6]),
  .ZN(_04369_)
);

NAND2_X1 _09951_ (
  .A1(_04368_),
  .A2(_04369_),
  .ZN(_04370_)
);

NAND2_X1 _09952_ (
  .A1(_04370_),
  .A2(_04338_),
  .ZN(_04371_)
);

NAND2_X1 _09953_ (
  .A1(_04351_),
  .A2(\sresult[55][6] ),
  .ZN(_04372_)
);

NAND2_X1 _09954_ (
  .A1(_04371_),
  .A2(_04372_),
  .ZN(_00666_)
);

NAND2_X1 _09955_ (
  .A1(_04346_),
  .A2(\sresult[54][7] ),
  .ZN(_04373_)
);

NAND2_X1 _09956_ (
  .A1(_04335_),
  .A2(din_21[7]),
  .ZN(_04374_)
);

NAND2_X1 _09957_ (
  .A1(_04373_),
  .A2(_04374_),
  .ZN(_04375_)
);

NAND2_X1 _09958_ (
  .A1(_04375_),
  .A2(_04338_),
  .ZN(_04376_)
);

NAND2_X1 _09959_ (
  .A1(_04351_),
  .A2(\sresult[55][7] ),
  .ZN(_04377_)
);

NAND2_X1 _09960_ (
  .A1(_04376_),
  .A2(_04377_),
  .ZN(_00667_)
);

NAND2_X1 _09961_ (
  .A1(_04346_),
  .A2(\sresult[54][8] ),
  .ZN(_04378_)
);

NAND2_X1 _09962_ (
  .A1(_04335_),
  .A2(din_21[8]),
  .ZN(_04379_)
);

NAND2_X1 _09963_ (
  .A1(_04378_),
  .A2(_04379_),
  .ZN(_04380_)
);

NAND2_X1 _09964_ (
  .A1(_04380_),
  .A2(_04338_),
  .ZN(_04381_)
);

NAND2_X1 _09965_ (
  .A1(_04351_),
  .A2(\sresult[55][8] ),
  .ZN(_04382_)
);

NAND2_X1 _09966_ (
  .A1(_04381_),
  .A2(_04382_),
  .ZN(_00668_)
);

NAND2_X1 _09967_ (
  .A1(_04346_),
  .A2(\sresult[54][9] ),
  .ZN(_04383_)
);

NAND2_X1 _09968_ (
  .A1(_04335_),
  .A2(din_21[9]),
  .ZN(_04384_)
);

NAND2_X1 _09969_ (
  .A1(_04383_),
  .A2(_04384_),
  .ZN(_04385_)
);

NAND2_X1 _09970_ (
  .A1(_04385_),
  .A2(_04338_),
  .ZN(_04386_)
);

NAND2_X1 _09971_ (
  .A1(_04351_),
  .A2(\sresult[55][9] ),
  .ZN(_04387_)
);

NAND2_X1 _09972_ (
  .A1(_04386_),
  .A2(_04387_),
  .ZN(_00669_)
);

NAND2_X1 _09973_ (
  .A1(_04346_),
  .A2(\sresult[54][10] ),
  .ZN(_04388_)
);

BUF_X4 _09974_ (
  .A(_04279_),
  .Z(_04389_)
);

NAND2_X1 _09975_ (
  .A1(_04389_),
  .A2(din_21[10]),
  .ZN(_04390_)
);

NAND2_X1 _09976_ (
  .A1(_04388_),
  .A2(_04390_),
  .ZN(_04391_)
);

BUF_X2 _09977_ (
  .A(_04172_),
  .Z(_04392_)
);

NAND2_X1 _09978_ (
  .A1(_04391_),
  .A2(_04392_),
  .ZN(_04393_)
);

NAND2_X1 _09979_ (
  .A1(_04351_),
  .A2(\sresult[55][10] ),
  .ZN(_04394_)
);

NAND2_X1 _09980_ (
  .A1(_04393_),
  .A2(_04394_),
  .ZN(_00670_)
);

NAND2_X1 _09981_ (
  .A1(_04346_),
  .A2(\sresult[54][11] ),
  .ZN(_04395_)
);

NAND2_X1 _09982_ (
  .A1(_04389_),
  .A2(din_21[11]),
  .ZN(_04396_)
);

NAND2_X1 _09983_ (
  .A1(_04395_),
  .A2(_04396_),
  .ZN(_04397_)
);

NAND2_X1 _09984_ (
  .A1(_04397_),
  .A2(_04392_),
  .ZN(_04398_)
);

NAND2_X1 _09985_ (
  .A1(_04351_),
  .A2(\sresult[55][11] ),
  .ZN(_04399_)
);

NAND2_X1 _09986_ (
  .A1(_04398_),
  .A2(_04399_),
  .ZN(_00671_)
);

BUF_X4 _09987_ (
  .A(_04235_),
  .Z(_04400_)
);

NAND2_X1 _09988_ (
  .A1(_04400_),
  .A2(\sresult[55][0] ),
  .ZN(_04401_)
);

NAND2_X1 _09989_ (
  .A1(_04389_),
  .A2(din_12[0]),
  .ZN(_04402_)
);

NAND2_X1 _09990_ (
  .A1(_04401_),
  .A2(_04402_),
  .ZN(_04403_)
);

NAND2_X1 _09991_ (
  .A1(_04403_),
  .A2(_04392_),
  .ZN(_04404_)
);

CLKBUF_X2 _09992_ (
  .A(_04296_),
  .Z(_04405_)
);

NAND2_X1 _09993_ (
  .A1(_04405_),
  .A2(\sresult[56][0] ),
  .ZN(_04406_)
);

NAND2_X1 _09994_ (
  .A1(_04404_),
  .A2(_04406_),
  .ZN(_00672_)
);

NAND2_X1 _09995_ (
  .A1(_04400_),
  .A2(\sresult[55][1] ),
  .ZN(_04407_)
);

NAND2_X1 _09996_ (
  .A1(_04389_),
  .A2(din_12[1]),
  .ZN(_04408_)
);

NAND2_X1 _09997_ (
  .A1(_04407_),
  .A2(_04408_),
  .ZN(_04409_)
);

NAND2_X1 _09998_ (
  .A1(_04409_),
  .A2(_04392_),
  .ZN(_04410_)
);

NAND2_X1 _09999_ (
  .A1(_04405_),
  .A2(\sresult[56][1] ),
  .ZN(_04411_)
);

NAND2_X1 _10000_ (
  .A1(_04410_),
  .A2(_04411_),
  .ZN(_00673_)
);

NAND2_X1 _10001_ (
  .A1(_04400_),
  .A2(\sresult[55][2] ),
  .ZN(_04412_)
);

NAND2_X1 _10002_ (
  .A1(_04389_),
  .A2(din_12[2]),
  .ZN(_04413_)
);

NAND2_X1 _10003_ (
  .A1(_04412_),
  .A2(_04413_),
  .ZN(_04414_)
);

NAND2_X1 _10004_ (
  .A1(_04414_),
  .A2(_04392_),
  .ZN(_04415_)
);

NAND2_X1 _10005_ (
  .A1(_04405_),
  .A2(\sresult[56][2] ),
  .ZN(_04416_)
);

NAND2_X1 _10006_ (
  .A1(_04415_),
  .A2(_04416_),
  .ZN(_00674_)
);

NAND2_X1 _10007_ (
  .A1(_04400_),
  .A2(\sresult[55][3] ),
  .ZN(_04417_)
);

NAND2_X1 _10008_ (
  .A1(_04389_),
  .A2(din_12[3]),
  .ZN(_04418_)
);

NAND2_X1 _10009_ (
  .A1(_04417_),
  .A2(_04418_),
  .ZN(_04419_)
);

NAND2_X1 _10010_ (
  .A1(_04419_),
  .A2(_04392_),
  .ZN(_04420_)
);

NAND2_X1 _10011_ (
  .A1(_04405_),
  .A2(\sresult[56][3] ),
  .ZN(_04421_)
);

NAND2_X1 _10012_ (
  .A1(_04420_),
  .A2(_04421_),
  .ZN(_00675_)
);

NAND2_X1 _10013_ (
  .A1(_04400_),
  .A2(\sresult[55][4] ),
  .ZN(_04422_)
);

NAND2_X1 _10014_ (
  .A1(_04389_),
  .A2(din_12[4]),
  .ZN(_04423_)
);

NAND2_X1 _10015_ (
  .A1(_04422_),
  .A2(_04423_),
  .ZN(_04424_)
);

NAND2_X1 _10016_ (
  .A1(_04424_),
  .A2(_04392_),
  .ZN(_04425_)
);

NAND2_X1 _10017_ (
  .A1(_04405_),
  .A2(\sresult[56][4] ),
  .ZN(_04426_)
);

NAND2_X1 _10018_ (
  .A1(_04425_),
  .A2(_04426_),
  .ZN(_00676_)
);

NAND2_X1 _10019_ (
  .A1(_04400_),
  .A2(\sresult[55][5] ),
  .ZN(_04427_)
);

NAND2_X1 _10020_ (
  .A1(_04389_),
  .A2(din_12[5]),
  .ZN(_04428_)
);

NAND2_X1 _10021_ (
  .A1(_04427_),
  .A2(_04428_),
  .ZN(_04429_)
);

NAND2_X1 _10022_ (
  .A1(_04429_),
  .A2(_04392_),
  .ZN(_04430_)
);

NAND2_X1 _10023_ (
  .A1(_04405_),
  .A2(\sresult[56][5] ),
  .ZN(_04431_)
);

NAND2_X1 _10024_ (
  .A1(_04430_),
  .A2(_04431_),
  .ZN(_00677_)
);

NAND2_X1 _10025_ (
  .A1(_04400_),
  .A2(\sresult[55][6] ),
  .ZN(_04432_)
);

NAND2_X1 _10026_ (
  .A1(_04389_),
  .A2(din_12[6]),
  .ZN(_04433_)
);

NAND2_X1 _10027_ (
  .A1(_04432_),
  .A2(_04433_),
  .ZN(_04434_)
);

NAND2_X1 _10028_ (
  .A1(_04434_),
  .A2(_04392_),
  .ZN(_04435_)
);

NAND2_X1 _10029_ (
  .A1(_04405_),
  .A2(\sresult[56][6] ),
  .ZN(_04436_)
);

NAND2_X1 _10030_ (
  .A1(_04435_),
  .A2(_04436_),
  .ZN(_00678_)
);

NAND2_X1 _10031_ (
  .A1(_04400_),
  .A2(\sresult[55][7] ),
  .ZN(_04437_)
);

NAND2_X1 _10032_ (
  .A1(_04389_),
  .A2(din_12[7]),
  .ZN(_04438_)
);

NAND2_X1 _10033_ (
  .A1(_04437_),
  .A2(_04438_),
  .ZN(_04439_)
);

NAND2_X1 _10034_ (
  .A1(_04439_),
  .A2(_04392_),
  .ZN(_04440_)
);

NAND2_X1 _10035_ (
  .A1(_04405_),
  .A2(\sresult[56][7] ),
  .ZN(_04441_)
);

NAND2_X1 _10036_ (
  .A1(_04440_),
  .A2(_04441_),
  .ZN(_00679_)
);

NAND2_X1 _10037_ (
  .A1(_04400_),
  .A2(\sresult[55][8] ),
  .ZN(_04442_)
);

BUF_X4 _10038_ (
  .A(_04279_),
  .Z(_04443_)
);

NAND2_X1 _10039_ (
  .A1(_04443_),
  .A2(din_12[8]),
  .ZN(_04444_)
);

NAND2_X1 _10040_ (
  .A1(_04442_),
  .A2(_04444_),
  .ZN(_04445_)
);

BUF_X2 _10041_ (
  .A(_04172_),
  .Z(_04446_)
);

NAND2_X1 _10042_ (
  .A1(_04445_),
  .A2(_04446_),
  .ZN(_04447_)
);

NAND2_X1 _10043_ (
  .A1(_04405_),
  .A2(\sresult[56][8] ),
  .ZN(_04448_)
);

NAND2_X1 _10044_ (
  .A1(_04447_),
  .A2(_04448_),
  .ZN(_00680_)
);

NAND2_X1 _10045_ (
  .A1(_04400_),
  .A2(\sresult[55][9] ),
  .ZN(_04449_)
);

NAND2_X1 _10046_ (
  .A1(_04443_),
  .A2(din_12[9]),
  .ZN(_04450_)
);

NAND2_X1 _10047_ (
  .A1(_04449_),
  .A2(_04450_),
  .ZN(_04451_)
);

NAND2_X1 _10048_ (
  .A1(_04451_),
  .A2(_04446_),
  .ZN(_04452_)
);

NAND2_X1 _10049_ (
  .A1(_04405_),
  .A2(\sresult[56][9] ),
  .ZN(_04453_)
);

NAND2_X1 _10050_ (
  .A1(_04452_),
  .A2(_04453_),
  .ZN(_00681_)
);

BUF_X4 _10051_ (
  .A(_04235_),
  .Z(_04454_)
);

NAND2_X1 _10052_ (
  .A1(_04454_),
  .A2(\sresult[55][10] ),
  .ZN(_04455_)
);

NAND2_X1 _10053_ (
  .A1(_04443_),
  .A2(din_12[10]),
  .ZN(_04456_)
);

NAND2_X1 _10054_ (
  .A1(_04455_),
  .A2(_04456_),
  .ZN(_04457_)
);

NAND2_X1 _10055_ (
  .A1(_04457_),
  .A2(_04446_),
  .ZN(_04458_)
);

CLKBUF_X2 _10056_ (
  .A(_04296_),
  .Z(_04459_)
);

NAND2_X1 _10057_ (
  .A1(_04459_),
  .A2(\sresult[56][10] ),
  .ZN(_04460_)
);

NAND2_X1 _10058_ (
  .A1(_04458_),
  .A2(_04460_),
  .ZN(_00682_)
);

NAND2_X1 _10059_ (
  .A1(_04454_),
  .A2(\sresult[55][11] ),
  .ZN(_04461_)
);

NAND2_X1 _10060_ (
  .A1(_04443_),
  .A2(din_12[11]),
  .ZN(_04462_)
);

NAND2_X1 _10061_ (
  .A1(_04461_),
  .A2(_04462_),
  .ZN(_04463_)
);

NAND2_X1 _10062_ (
  .A1(_04463_),
  .A2(_04446_),
  .ZN(_04464_)
);

NAND2_X1 _10063_ (
  .A1(_04459_),
  .A2(\sresult[56][11] ),
  .ZN(_04465_)
);

NAND2_X1 _10064_ (
  .A1(_04464_),
  .A2(_04465_),
  .ZN(_00683_)
);

NAND2_X1 _10065_ (
  .A1(_04454_),
  .A2(\sresult[56][0] ),
  .ZN(_04466_)
);

NAND2_X1 _10066_ (
  .A1(_04443_),
  .A2(din_03[0]),
  .ZN(_04467_)
);

NAND2_X1 _10067_ (
  .A1(_04466_),
  .A2(_04467_),
  .ZN(_04468_)
);

NAND2_X1 _10068_ (
  .A1(_04468_),
  .A2(_04446_),
  .ZN(_04469_)
);

NAND2_X1 _10069_ (
  .A1(_04459_),
  .A2(\sresult[57][0] ),
  .ZN(_04470_)
);

NAND2_X1 _10070_ (
  .A1(_04469_),
  .A2(_04470_),
  .ZN(_00684_)
);

NAND2_X1 _10071_ (
  .A1(_04454_),
  .A2(\sresult[56][1] ),
  .ZN(_04471_)
);

NAND2_X1 _10072_ (
  .A1(_04443_),
  .A2(din_03[1]),
  .ZN(_04472_)
);

NAND2_X1 _10073_ (
  .A1(_04471_),
  .A2(_04472_),
  .ZN(_04473_)
);

NAND2_X1 _10074_ (
  .A1(_04473_),
  .A2(_04446_),
  .ZN(_04474_)
);

NAND2_X1 _10075_ (
  .A1(_04459_),
  .A2(\sresult[57][1] ),
  .ZN(_04475_)
);

NAND2_X1 _10076_ (
  .A1(_04474_),
  .A2(_04475_),
  .ZN(_00685_)
);

NAND2_X1 _10077_ (
  .A1(_04454_),
  .A2(\sresult[56][2] ),
  .ZN(_04476_)
);

NAND2_X1 _10078_ (
  .A1(_04443_),
  .A2(din_03[2]),
  .ZN(_04477_)
);

NAND2_X1 _10079_ (
  .A1(_04476_),
  .A2(_04477_),
  .ZN(_04478_)
);

NAND2_X1 _10080_ (
  .A1(_04478_),
  .A2(_04446_),
  .ZN(_04479_)
);

NAND2_X1 _10081_ (
  .A1(_04459_),
  .A2(\sresult[57][2] ),
  .ZN(_04480_)
);

NAND2_X1 _10082_ (
  .A1(_04479_),
  .A2(_04480_),
  .ZN(_00686_)
);

NAND2_X1 _10083_ (
  .A1(_04454_),
  .A2(\sresult[56][3] ),
  .ZN(_04481_)
);

NAND2_X1 _10084_ (
  .A1(_04443_),
  .A2(din_03[3]),
  .ZN(_04482_)
);

NAND2_X1 _10085_ (
  .A1(_04481_),
  .A2(_04482_),
  .ZN(_04483_)
);

NAND2_X1 _10086_ (
  .A1(_04483_),
  .A2(_04446_),
  .ZN(_04484_)
);

NAND2_X1 _10087_ (
  .A1(_04459_),
  .A2(\sresult[57][3] ),
  .ZN(_04485_)
);

NAND2_X1 _10088_ (
  .A1(_04484_),
  .A2(_04485_),
  .ZN(_00687_)
);

NAND2_X1 _10089_ (
  .A1(_04454_),
  .A2(\sresult[56][4] ),
  .ZN(_04486_)
);

NAND2_X1 _10090_ (
  .A1(_04443_),
  .A2(din_03[4]),
  .ZN(_04487_)
);

NAND2_X1 _10091_ (
  .A1(_04486_),
  .A2(_04487_),
  .ZN(_04488_)
);

NAND2_X1 _10092_ (
  .A1(_04488_),
  .A2(_04446_),
  .ZN(_04489_)
);

NAND2_X1 _10093_ (
  .A1(_04459_),
  .A2(\sresult[57][4] ),
  .ZN(_04490_)
);

NAND2_X1 _10094_ (
  .A1(_04489_),
  .A2(_04490_),
  .ZN(_00688_)
);

NAND2_X1 _10095_ (
  .A1(_04454_),
  .A2(\sresult[56][5] ),
  .ZN(_04491_)
);

NAND2_X1 _10096_ (
  .A1(_04443_),
  .A2(din_03[5]),
  .ZN(_04492_)
);

NAND2_X1 _10097_ (
  .A1(_04491_),
  .A2(_04492_),
  .ZN(_04493_)
);

NAND2_X1 _10098_ (
  .A1(_04493_),
  .A2(_04446_),
  .ZN(_04494_)
);

NAND2_X1 _10099_ (
  .A1(_04459_),
  .A2(\sresult[57][5] ),
  .ZN(_04495_)
);

NAND2_X1 _10100_ (
  .A1(_04494_),
  .A2(_04495_),
  .ZN(_00689_)
);

NAND2_X1 _10101_ (
  .A1(_04454_),
  .A2(\sresult[56][6] ),
  .ZN(_04496_)
);

BUF_X4 _10102_ (
  .A(_04279_),
  .Z(_04497_)
);

NAND2_X1 _10103_ (
  .A1(_04497_),
  .A2(din_03[6]),
  .ZN(_04498_)
);

NAND2_X1 _10104_ (
  .A1(_04496_),
  .A2(_04498_),
  .ZN(_04499_)
);

BUF_X2 _10105_ (
  .A(_04172_),
  .Z(_04500_)
);

NAND2_X1 _10106_ (
  .A1(_04499_),
  .A2(_04500_),
  .ZN(_04501_)
);

NAND2_X1 _10107_ (
  .A1(_04459_),
  .A2(\sresult[57][6] ),
  .ZN(_04502_)
);

NAND2_X1 _10108_ (
  .A1(_04501_),
  .A2(_04502_),
  .ZN(_00690_)
);

NAND2_X1 _10109_ (
  .A1(_04454_),
  .A2(\sresult[56][7] ),
  .ZN(_04503_)
);

NAND2_X1 _10110_ (
  .A1(_04497_),
  .A2(din_03[7]),
  .ZN(_04504_)
);

NAND2_X1 _10111_ (
  .A1(_04503_),
  .A2(_04504_),
  .ZN(_04505_)
);

NAND2_X1 _10112_ (
  .A1(_04505_),
  .A2(_04500_),
  .ZN(_04506_)
);

NAND2_X1 _10113_ (
  .A1(_04459_),
  .A2(\sresult[57][7] ),
  .ZN(_04507_)
);

NAND2_X1 _10114_ (
  .A1(_04506_),
  .A2(_04507_),
  .ZN(_00691_)
);

BUF_X4 _10115_ (
  .A(_04235_),
  .Z(_04508_)
);

NAND2_X1 _10116_ (
  .A1(_04508_),
  .A2(\sresult[56][8] ),
  .ZN(_04509_)
);

NAND2_X1 _10117_ (
  .A1(_04497_),
  .A2(din_03[8]),
  .ZN(_04510_)
);

NAND2_X1 _10118_ (
  .A1(_04509_),
  .A2(_04510_),
  .ZN(_04511_)
);

NAND2_X1 _10119_ (
  .A1(_04511_),
  .A2(_04500_),
  .ZN(_04512_)
);

CLKBUF_X2 _10120_ (
  .A(_04296_),
  .Z(_04513_)
);

NAND2_X1 _10121_ (
  .A1(_04513_),
  .A2(\sresult[57][8] ),
  .ZN(_04514_)
);

NAND2_X1 _10122_ (
  .A1(_04512_),
  .A2(_04514_),
  .ZN(_00692_)
);

NAND2_X1 _10123_ (
  .A1(_04508_),
  .A2(\sresult[56][9] ),
  .ZN(_04515_)
);

NAND2_X1 _10124_ (
  .A1(_04497_),
  .A2(din_03[9]),
  .ZN(_04516_)
);

NAND2_X1 _10125_ (
  .A1(_04515_),
  .A2(_04516_),
  .ZN(_04517_)
);

NAND2_X1 _10126_ (
  .A1(_04517_),
  .A2(_04500_),
  .ZN(_04518_)
);

NAND2_X1 _10127_ (
  .A1(_04513_),
  .A2(\sresult[57][9] ),
  .ZN(_04519_)
);

NAND2_X1 _10128_ (
  .A1(_04518_),
  .A2(_04519_),
  .ZN(_00693_)
);

NAND2_X1 _10129_ (
  .A1(_04508_),
  .A2(\sresult[56][10] ),
  .ZN(_04520_)
);

NAND2_X1 _10130_ (
  .A1(_04497_),
  .A2(din_03[10]),
  .ZN(_04521_)
);

NAND2_X1 _10131_ (
  .A1(_04520_),
  .A2(_04521_),
  .ZN(_04522_)
);

NAND2_X1 _10132_ (
  .A1(_04522_),
  .A2(_04500_),
  .ZN(_04523_)
);

NAND2_X1 _10133_ (
  .A1(_04513_),
  .A2(\sresult[57][10] ),
  .ZN(_04524_)
);

NAND2_X1 _10134_ (
  .A1(_04523_),
  .A2(_04524_),
  .ZN(_00694_)
);

NAND2_X1 _10135_ (
  .A1(_04508_),
  .A2(\sresult[56][11] ),
  .ZN(_04525_)
);

NAND2_X1 _10136_ (
  .A1(_04497_),
  .A2(din_03[11]),
  .ZN(_04526_)
);

NAND2_X1 _10137_ (
  .A1(_04525_),
  .A2(_04526_),
  .ZN(_04527_)
);

NAND2_X1 _10138_ (
  .A1(_04527_),
  .A2(_04500_),
  .ZN(_04528_)
);

NAND2_X1 _10139_ (
  .A1(_04513_),
  .A2(\sresult[57][11] ),
  .ZN(_04529_)
);

NAND2_X1 _10140_ (
  .A1(_04528_),
  .A2(_04529_),
  .ZN(_00695_)
);

NAND2_X1 _10141_ (
  .A1(_04508_),
  .A2(\sresult[57][0] ),
  .ZN(_04530_)
);

NAND2_X1 _10142_ (
  .A1(_04497_),
  .A2(din_02[0]),
  .ZN(_04531_)
);

NAND2_X1 _10143_ (
  .A1(_04530_),
  .A2(_04531_),
  .ZN(_04532_)
);

NAND2_X1 _10144_ (
  .A1(_04532_),
  .A2(_04500_),
  .ZN(_04533_)
);

NAND2_X1 _10145_ (
  .A1(_04513_),
  .A2(\sresult[58][0] ),
  .ZN(_04534_)
);

NAND2_X1 _10146_ (
  .A1(_04533_),
  .A2(_04534_),
  .ZN(_00696_)
);

NAND2_X1 _10147_ (
  .A1(_04508_),
  .A2(\sresult[57][1] ),
  .ZN(_04535_)
);

NAND2_X1 _10148_ (
  .A1(_04497_),
  .A2(din_02[1]),
  .ZN(_04536_)
);

NAND2_X1 _10149_ (
  .A1(_04535_),
  .A2(_04536_),
  .ZN(_04537_)
);

NAND2_X1 _10150_ (
  .A1(_04537_),
  .A2(_04500_),
  .ZN(_04538_)
);

NAND2_X1 _10151_ (
  .A1(_04513_),
  .A2(\sresult[58][1] ),
  .ZN(_04539_)
);

NAND2_X1 _10152_ (
  .A1(_04538_),
  .A2(_04539_),
  .ZN(_00697_)
);

NAND2_X1 _10153_ (
  .A1(_04508_),
  .A2(\sresult[57][2] ),
  .ZN(_04540_)
);

NAND2_X1 _10154_ (
  .A1(_04497_),
  .A2(din_02[2]),
  .ZN(_04541_)
);

NAND2_X1 _10155_ (
  .A1(_04540_),
  .A2(_04541_),
  .ZN(_04542_)
);

NAND2_X1 _10156_ (
  .A1(_04542_),
  .A2(_04500_),
  .ZN(_04543_)
);

NAND2_X1 _10157_ (
  .A1(_04513_),
  .A2(\sresult[58][2] ),
  .ZN(_04544_)
);

NAND2_X1 _10158_ (
  .A1(_04543_),
  .A2(_04544_),
  .ZN(_00698_)
);

NAND2_X1 _10159_ (
  .A1(_04508_),
  .A2(\sresult[57][3] ),
  .ZN(_04545_)
);

NAND2_X1 _10160_ (
  .A1(_04497_),
  .A2(din_02[3]),
  .ZN(_04546_)
);

NAND2_X1 _10161_ (
  .A1(_04545_),
  .A2(_04546_),
  .ZN(_04547_)
);

NAND2_X1 _10162_ (
  .A1(_04547_),
  .A2(_04500_),
  .ZN(_04548_)
);

NAND2_X1 _10163_ (
  .A1(_04513_),
  .A2(\sresult[58][3] ),
  .ZN(_04549_)
);

NAND2_X1 _10164_ (
  .A1(_04548_),
  .A2(_04549_),
  .ZN(_00699_)
);

NAND2_X1 _10165_ (
  .A1(_04508_),
  .A2(\sresult[57][4] ),
  .ZN(_04550_)
);

BUF_X4 _10166_ (
  .A(_04279_),
  .Z(_04551_)
);

NAND2_X1 _10167_ (
  .A1(_04551_),
  .A2(din_02[4]),
  .ZN(_04552_)
);

NAND2_X1 _10168_ (
  .A1(_04550_),
  .A2(_04552_),
  .ZN(_04553_)
);

BUF_X2 _10169_ (
  .A(_04172_),
  .Z(_04554_)
);

NAND2_X1 _10170_ (
  .A1(_04553_),
  .A2(_04554_),
  .ZN(_04555_)
);

NAND2_X1 _10171_ (
  .A1(_04513_),
  .A2(\sresult[58][4] ),
  .ZN(_04556_)
);

NAND2_X1 _10172_ (
  .A1(_04555_),
  .A2(_04556_),
  .ZN(_00700_)
);

NAND2_X1 _10173_ (
  .A1(_04508_),
  .A2(\sresult[57][5] ),
  .ZN(_04557_)
);

NAND2_X1 _10174_ (
  .A1(_04551_),
  .A2(din_02[5]),
  .ZN(_04558_)
);

NAND2_X1 _10175_ (
  .A1(_04557_),
  .A2(_04558_),
  .ZN(_04559_)
);

NAND2_X1 _10176_ (
  .A1(_04559_),
  .A2(_04554_),
  .ZN(_04560_)
);

NAND2_X1 _10177_ (
  .A1(_04513_),
  .A2(\sresult[58][5] ),
  .ZN(_04561_)
);

NAND2_X1 _10178_ (
  .A1(_04560_),
  .A2(_04561_),
  .ZN(_00701_)
);

BUF_X4 _10179_ (
  .A(_04235_),
  .Z(_04562_)
);

NAND2_X1 _10180_ (
  .A1(_04562_),
  .A2(\sresult[57][6] ),
  .ZN(_04563_)
);

NAND2_X1 _10181_ (
  .A1(_04551_),
  .A2(din_02[6]),
  .ZN(_04564_)
);

NAND2_X1 _10182_ (
  .A1(_04563_),
  .A2(_04564_),
  .ZN(_04565_)
);

NAND2_X1 _10183_ (
  .A1(_04565_),
  .A2(_04554_),
  .ZN(_04566_)
);

CLKBUF_X2 _10184_ (
  .A(_04296_),
  .Z(_04567_)
);

NAND2_X1 _10185_ (
  .A1(_04567_),
  .A2(\sresult[58][6] ),
  .ZN(_04568_)
);

NAND2_X1 _10186_ (
  .A1(_04566_),
  .A2(_04568_),
  .ZN(_00702_)
);

NAND2_X1 _10187_ (
  .A1(_04562_),
  .A2(\sresult[57][7] ),
  .ZN(_04569_)
);

NAND2_X1 _10188_ (
  .A1(_04551_),
  .A2(din_02[7]),
  .ZN(_04570_)
);

NAND2_X1 _10189_ (
  .A1(_04569_),
  .A2(_04570_),
  .ZN(_04571_)
);

NAND2_X1 _10190_ (
  .A1(_04571_),
  .A2(_04554_),
  .ZN(_04572_)
);

NAND2_X1 _10191_ (
  .A1(_04567_),
  .A2(\sresult[58][7] ),
  .ZN(_04573_)
);

NAND2_X1 _10192_ (
  .A1(_04572_),
  .A2(_04573_),
  .ZN(_00703_)
);

NAND2_X1 _10193_ (
  .A1(_04562_),
  .A2(\sresult[57][8] ),
  .ZN(_04574_)
);

NAND2_X1 _10194_ (
  .A1(_04551_),
  .A2(din_02[8]),
  .ZN(_04575_)
);

NAND2_X1 _10195_ (
  .A1(_04574_),
  .A2(_04575_),
  .ZN(_04576_)
);

NAND2_X1 _10196_ (
  .A1(_04576_),
  .A2(_04554_),
  .ZN(_04577_)
);

NAND2_X1 _10197_ (
  .A1(_04567_),
  .A2(\sresult[58][8] ),
  .ZN(_04578_)
);

NAND2_X1 _10198_ (
  .A1(_04577_),
  .A2(_04578_),
  .ZN(_00704_)
);

NAND2_X1 _10199_ (
  .A1(_04562_),
  .A2(\sresult[57][9] ),
  .ZN(_04579_)
);

NAND2_X1 _10200_ (
  .A1(_04551_),
  .A2(din_02[9]),
  .ZN(_04580_)
);

NAND2_X1 _10201_ (
  .A1(_04579_),
  .A2(_04580_),
  .ZN(_04581_)
);

NAND2_X1 _10202_ (
  .A1(_04581_),
  .A2(_04554_),
  .ZN(_04582_)
);

NAND2_X1 _10203_ (
  .A1(_04567_),
  .A2(\sresult[58][9] ),
  .ZN(_04583_)
);

NAND2_X1 _10204_ (
  .A1(_04582_),
  .A2(_04583_),
  .ZN(_00705_)
);

NAND2_X1 _10205_ (
  .A1(_04562_),
  .A2(\sresult[57][10] ),
  .ZN(_04584_)
);

NAND2_X1 _10206_ (
  .A1(_04551_),
  .A2(din_02[10]),
  .ZN(_04585_)
);

NAND2_X1 _10207_ (
  .A1(_04584_),
  .A2(_04585_),
  .ZN(_04586_)
);

NAND2_X1 _10208_ (
  .A1(_04586_),
  .A2(_04554_),
  .ZN(_04587_)
);

NAND2_X1 _10209_ (
  .A1(_04567_),
  .A2(\sresult[58][10] ),
  .ZN(_04588_)
);

NAND2_X1 _10210_ (
  .A1(_04587_),
  .A2(_04588_),
  .ZN(_00706_)
);

NAND2_X1 _10211_ (
  .A1(_04562_),
  .A2(\sresult[57][11] ),
  .ZN(_04589_)
);

NAND2_X1 _10212_ (
  .A1(_04551_),
  .A2(din_02[11]),
  .ZN(_04590_)
);

NAND2_X1 _10213_ (
  .A1(_04589_),
  .A2(_04590_),
  .ZN(_04591_)
);

NAND2_X1 _10214_ (
  .A1(_04591_),
  .A2(_04554_),
  .ZN(_04592_)
);

NAND2_X1 _10215_ (
  .A1(_04567_),
  .A2(\sresult[58][11] ),
  .ZN(_04593_)
);

NAND2_X1 _10216_ (
  .A1(_04592_),
  .A2(_04593_),
  .ZN(_00707_)
);

NAND2_X1 _10217_ (
  .A1(_04562_),
  .A2(\sresult[58][0] ),
  .ZN(_04594_)
);

NAND2_X1 _10218_ (
  .A1(_04551_),
  .A2(din_11[0]),
  .ZN(_04595_)
);

NAND2_X1 _10219_ (
  .A1(_04594_),
  .A2(_04595_),
  .ZN(_04596_)
);

NAND2_X1 _10220_ (
  .A1(_04596_),
  .A2(_04554_),
  .ZN(_04597_)
);

NAND2_X1 _10221_ (
  .A1(_04567_),
  .A2(\sresult[59][0] ),
  .ZN(_04598_)
);

NAND2_X1 _10222_ (
  .A1(_04597_),
  .A2(_04598_),
  .ZN(_00708_)
);

NAND2_X1 _10223_ (
  .A1(_04562_),
  .A2(\sresult[58][1] ),
  .ZN(_04599_)
);

NAND2_X1 _10224_ (
  .A1(_04551_),
  .A2(din_11[1]),
  .ZN(_04600_)
);

NAND2_X1 _10225_ (
  .A1(_04599_),
  .A2(_04600_),
  .ZN(_04601_)
);

NAND2_X1 _10226_ (
  .A1(_04601_),
  .A2(_04554_),
  .ZN(_04602_)
);

NAND2_X1 _10227_ (
  .A1(_04567_),
  .A2(\sresult[59][1] ),
  .ZN(_04603_)
);

NAND2_X1 _10228_ (
  .A1(_04602_),
  .A2(_04603_),
  .ZN(_00709_)
);

NAND2_X1 _10229_ (
  .A1(_04562_),
  .A2(\sresult[58][2] ),
  .ZN(_04604_)
);

BUF_X4 _10230_ (
  .A(_04279_),
  .Z(_04605_)
);

NAND2_X1 _10231_ (
  .A1(_04605_),
  .A2(din_11[2]),
  .ZN(_04606_)
);

NAND2_X1 _10232_ (
  .A1(_04604_),
  .A2(_04606_),
  .ZN(_04607_)
);

BUF_X2 _10233_ (
  .A(_04172_),
  .Z(_04608_)
);

NAND2_X1 _10234_ (
  .A1(_04607_),
  .A2(_04608_),
  .ZN(_04609_)
);

NAND2_X1 _10235_ (
  .A1(_04567_),
  .A2(\sresult[59][2] ),
  .ZN(_04610_)
);

NAND2_X1 _10236_ (
  .A1(_04609_),
  .A2(_04610_),
  .ZN(_00710_)
);

NAND2_X1 _10237_ (
  .A1(_04562_),
  .A2(\sresult[58][3] ),
  .ZN(_04611_)
);

NAND2_X1 _10238_ (
  .A1(_04605_),
  .A2(din_11[3]),
  .ZN(_04612_)
);

NAND2_X1 _10239_ (
  .A1(_04611_),
  .A2(_04612_),
  .ZN(_04613_)
);

NAND2_X1 _10240_ (
  .A1(_04613_),
  .A2(_04608_),
  .ZN(_04614_)
);

NAND2_X1 _10241_ (
  .A1(_04567_),
  .A2(\sresult[59][3] ),
  .ZN(_04615_)
);

NAND2_X1 _10242_ (
  .A1(_04614_),
  .A2(_04615_),
  .ZN(_00711_)
);

BUF_X4 _10243_ (
  .A(_04235_),
  .Z(_04616_)
);

NAND2_X1 _10244_ (
  .A1(_04616_),
  .A2(\sresult[58][4] ),
  .ZN(_04617_)
);

NAND2_X1 _10245_ (
  .A1(_04605_),
  .A2(din_11[4]),
  .ZN(_04618_)
);

NAND2_X1 _10246_ (
  .A1(_04617_),
  .A2(_04618_),
  .ZN(_04619_)
);

NAND2_X1 _10247_ (
  .A1(_04619_),
  .A2(_04608_),
  .ZN(_04620_)
);

CLKBUF_X2 _10248_ (
  .A(_04296_),
  .Z(_04621_)
);

NAND2_X1 _10249_ (
  .A1(_04621_),
  .A2(\sresult[59][4] ),
  .ZN(_04622_)
);

NAND2_X1 _10250_ (
  .A1(_04620_),
  .A2(_04622_),
  .ZN(_00712_)
);

NAND2_X1 _10251_ (
  .A1(_04616_),
  .A2(\sresult[58][5] ),
  .ZN(_04623_)
);

NAND2_X1 _10252_ (
  .A1(_04605_),
  .A2(din_11[5]),
  .ZN(_04624_)
);

NAND2_X1 _10253_ (
  .A1(_04623_),
  .A2(_04624_),
  .ZN(_04625_)
);

NAND2_X1 _10254_ (
  .A1(_04625_),
  .A2(_04608_),
  .ZN(_04626_)
);

NAND2_X1 _10255_ (
  .A1(_04621_),
  .A2(\sresult[59][5] ),
  .ZN(_04627_)
);

NAND2_X1 _10256_ (
  .A1(_04626_),
  .A2(_04627_),
  .ZN(_00713_)
);

NAND2_X1 _10257_ (
  .A1(_04616_),
  .A2(\sresult[58][6] ),
  .ZN(_04628_)
);

NAND2_X1 _10258_ (
  .A1(_04605_),
  .A2(din_11[6]),
  .ZN(_04629_)
);

NAND2_X1 _10259_ (
  .A1(_04628_),
  .A2(_04629_),
  .ZN(_04630_)
);

NAND2_X1 _10260_ (
  .A1(_04630_),
  .A2(_04608_),
  .ZN(_04631_)
);

NAND2_X1 _10261_ (
  .A1(_04621_),
  .A2(\sresult[59][6] ),
  .ZN(_04632_)
);

NAND2_X1 _10262_ (
  .A1(_04631_),
  .A2(_04632_),
  .ZN(_00714_)
);

NAND2_X1 _10263_ (
  .A1(_04616_),
  .A2(\sresult[58][7] ),
  .ZN(_04633_)
);

NAND2_X1 _10264_ (
  .A1(_04605_),
  .A2(din_11[7]),
  .ZN(_04634_)
);

NAND2_X1 _10265_ (
  .A1(_04633_),
  .A2(_04634_),
  .ZN(_04635_)
);

NAND2_X1 _10266_ (
  .A1(_04635_),
  .A2(_04608_),
  .ZN(_04636_)
);

NAND2_X1 _10267_ (
  .A1(_04621_),
  .A2(\sresult[59][7] ),
  .ZN(_04637_)
);

NAND2_X1 _10268_ (
  .A1(_04636_),
  .A2(_04637_),
  .ZN(_00715_)
);

NAND2_X1 _10269_ (
  .A1(_04616_),
  .A2(\sresult[58][8] ),
  .ZN(_04638_)
);

NAND2_X1 _10270_ (
  .A1(_04605_),
  .A2(din_11[8]),
  .ZN(_04639_)
);

NAND2_X1 _10271_ (
  .A1(_04638_),
  .A2(_04639_),
  .ZN(_04640_)
);

NAND2_X1 _10272_ (
  .A1(_04640_),
  .A2(_04608_),
  .ZN(_04641_)
);

NAND2_X1 _10273_ (
  .A1(_04621_),
  .A2(\sresult[59][8] ),
  .ZN(_04642_)
);

NAND2_X1 _10274_ (
  .A1(_04641_),
  .A2(_04642_),
  .ZN(_00716_)
);

NAND2_X1 _10275_ (
  .A1(_04616_),
  .A2(\sresult[58][9] ),
  .ZN(_04643_)
);

NAND2_X1 _10276_ (
  .A1(_04605_),
  .A2(din_11[9]),
  .ZN(_04644_)
);

NAND2_X1 _10277_ (
  .A1(_04643_),
  .A2(_04644_),
  .ZN(_04645_)
);

NAND2_X1 _10278_ (
  .A1(_04645_),
  .A2(_04608_),
  .ZN(_04646_)
);

NAND2_X1 _10279_ (
  .A1(_04621_),
  .A2(\sresult[59][9] ),
  .ZN(_04647_)
);

NAND2_X1 _10280_ (
  .A1(_04646_),
  .A2(_04647_),
  .ZN(_00717_)
);

NAND2_X1 _10281_ (
  .A1(_04616_),
  .A2(\sresult[58][10] ),
  .ZN(_04648_)
);

NAND2_X1 _10282_ (
  .A1(_04605_),
  .A2(din_11[10]),
  .ZN(_04649_)
);

NAND2_X1 _10283_ (
  .A1(_04648_),
  .A2(_04649_),
  .ZN(_04650_)
);

NAND2_X1 _10284_ (
  .A1(_04650_),
  .A2(_04608_),
  .ZN(_04651_)
);

NAND2_X1 _10285_ (
  .A1(_04621_),
  .A2(\sresult[59][10] ),
  .ZN(_04652_)
);

NAND2_X1 _10286_ (
  .A1(_04651_),
  .A2(_04652_),
  .ZN(_00718_)
);

NAND2_X1 _10287_ (
  .A1(_04616_),
  .A2(\sresult[58][11] ),
  .ZN(_04653_)
);

NAND2_X1 _10288_ (
  .A1(_04605_),
  .A2(din_11[11]),
  .ZN(_04654_)
);

NAND2_X1 _10289_ (
  .A1(_04653_),
  .A2(_04654_),
  .ZN(_04655_)
);

NAND2_X1 _10290_ (
  .A1(_04655_),
  .A2(_04608_),
  .ZN(_04656_)
);

NAND2_X1 _10291_ (
  .A1(_04621_),
  .A2(\sresult[59][11] ),
  .ZN(_04657_)
);

NAND2_X1 _10292_ (
  .A1(_04656_),
  .A2(_04657_),
  .ZN(_00719_)
);

NAND2_X1 _10293_ (
  .A1(_04616_),
  .A2(\sresult[59][0] ),
  .ZN(_04658_)
);

BUF_X4 _10294_ (
  .A(_04279_),
  .Z(_04659_)
);

NAND2_X1 _10295_ (
  .A1(_04659_),
  .A2(din_20[0]),
  .ZN(_04660_)
);

NAND2_X1 _10296_ (
  .A1(_04658_),
  .A2(_04660_),
  .ZN(_04661_)
);

BUF_X2 _10297_ (
  .A(_04172_),
  .Z(_04662_)
);

NAND2_X1 _10298_ (
  .A1(_04661_),
  .A2(_04662_),
  .ZN(_04663_)
);

NAND2_X1 _10299_ (
  .A1(_04621_),
  .A2(\sresult[60][0] ),
  .ZN(_04664_)
);

NAND2_X1 _10300_ (
  .A1(_04663_),
  .A2(_04664_),
  .ZN(_00720_)
);

NAND2_X1 _10301_ (
  .A1(_04616_),
  .A2(\sresult[59][1] ),
  .ZN(_04665_)
);

NAND2_X1 _10302_ (
  .A1(_04659_),
  .A2(din_20[1]),
  .ZN(_04666_)
);

NAND2_X1 _10303_ (
  .A1(_04665_),
  .A2(_04666_),
  .ZN(_04667_)
);

NAND2_X1 _10304_ (
  .A1(_04667_),
  .A2(_04662_),
  .ZN(_04668_)
);

NAND2_X1 _10305_ (
  .A1(_04621_),
  .A2(\sresult[60][1] ),
  .ZN(_04669_)
);

NAND2_X1 _10306_ (
  .A1(_04668_),
  .A2(_04669_),
  .ZN(_00721_)
);

BUF_X4 _10307_ (
  .A(_04235_),
  .Z(_04670_)
);

NAND2_X1 _10308_ (
  .A1(_04670_),
  .A2(\sresult[59][2] ),
  .ZN(_04671_)
);

NAND2_X1 _10309_ (
  .A1(_04659_),
  .A2(din_20[2]),
  .ZN(_04672_)
);

NAND2_X1 _10310_ (
  .A1(_04671_),
  .A2(_04672_),
  .ZN(_04673_)
);

NAND2_X1 _10311_ (
  .A1(_04673_),
  .A2(_04662_),
  .ZN(_04674_)
);

CLKBUF_X2 _10312_ (
  .A(_04296_),
  .Z(_04675_)
);

NAND2_X1 _10313_ (
  .A1(_04675_),
  .A2(\sresult[60][2] ),
  .ZN(_04676_)
);

NAND2_X1 _10314_ (
  .A1(_04674_),
  .A2(_04676_),
  .ZN(_00722_)
);

NAND2_X1 _10315_ (
  .A1(_04670_),
  .A2(\sresult[59][3] ),
  .ZN(_04677_)
);

NAND2_X1 _10316_ (
  .A1(_04659_),
  .A2(din_20[3]),
  .ZN(_04678_)
);

NAND2_X1 _10317_ (
  .A1(_04677_),
  .A2(_04678_),
  .ZN(_04679_)
);

NAND2_X1 _10318_ (
  .A1(_04679_),
  .A2(_04662_),
  .ZN(_04680_)
);

NAND2_X1 _10319_ (
  .A1(_04675_),
  .A2(\sresult[60][3] ),
  .ZN(_04681_)
);

NAND2_X1 _10320_ (
  .A1(_04680_),
  .A2(_04681_),
  .ZN(_00723_)
);

NAND2_X1 _10321_ (
  .A1(_04670_),
  .A2(\sresult[59][4] ),
  .ZN(_04682_)
);

NAND2_X1 _10322_ (
  .A1(_04659_),
  .A2(din_20[4]),
  .ZN(_04683_)
);

NAND2_X1 _10323_ (
  .A1(_04682_),
  .A2(_04683_),
  .ZN(_04684_)
);

NAND2_X1 _10324_ (
  .A1(_04684_),
  .A2(_04662_),
  .ZN(_04685_)
);

NAND2_X1 _10325_ (
  .A1(_04675_),
  .A2(\sresult[60][4] ),
  .ZN(_04686_)
);

NAND2_X1 _10326_ (
  .A1(_04685_),
  .A2(_04686_),
  .ZN(_00724_)
);

NAND2_X1 _10327_ (
  .A1(_04670_),
  .A2(\sresult[59][5] ),
  .ZN(_04687_)
);

NAND2_X1 _10328_ (
  .A1(_04659_),
  .A2(din_20[5]),
  .ZN(_04688_)
);

NAND2_X1 _10329_ (
  .A1(_04687_),
  .A2(_04688_),
  .ZN(_04689_)
);

NAND2_X1 _10330_ (
  .A1(_04689_),
  .A2(_04662_),
  .ZN(_04690_)
);

NAND2_X1 _10331_ (
  .A1(_04675_),
  .A2(\sresult[60][5] ),
  .ZN(_04691_)
);

NAND2_X1 _10332_ (
  .A1(_04690_),
  .A2(_04691_),
  .ZN(_00725_)
);

NAND2_X1 _10333_ (
  .A1(_04670_),
  .A2(\sresult[59][6] ),
  .ZN(_04692_)
);

NAND2_X1 _10334_ (
  .A1(_04659_),
  .A2(din_20[6]),
  .ZN(_04693_)
);

NAND2_X1 _10335_ (
  .A1(_04692_),
  .A2(_04693_),
  .ZN(_04694_)
);

NAND2_X1 _10336_ (
  .A1(_04694_),
  .A2(_04662_),
  .ZN(_04695_)
);

NAND2_X1 _10337_ (
  .A1(_04675_),
  .A2(\sresult[60][6] ),
  .ZN(_04696_)
);

NAND2_X1 _10338_ (
  .A1(_04695_),
  .A2(_04696_),
  .ZN(_00726_)
);

NAND2_X1 _10339_ (
  .A1(_04670_),
  .A2(\sresult[59][7] ),
  .ZN(_04697_)
);

NAND2_X1 _10340_ (
  .A1(_04659_),
  .A2(din_20[7]),
  .ZN(_04698_)
);

NAND2_X1 _10341_ (
  .A1(_04697_),
  .A2(_04698_),
  .ZN(_04699_)
);

NAND2_X1 _10342_ (
  .A1(_04699_),
  .A2(_04662_),
  .ZN(_04700_)
);

NAND2_X1 _10343_ (
  .A1(_04675_),
  .A2(\sresult[60][7] ),
  .ZN(_04701_)
);

NAND2_X1 _10344_ (
  .A1(_04700_),
  .A2(_04701_),
  .ZN(_00727_)
);

NAND2_X1 _10345_ (
  .A1(_04670_),
  .A2(\sresult[59][8] ),
  .ZN(_04702_)
);

NAND2_X1 _10346_ (
  .A1(_04659_),
  .A2(din_20[8]),
  .ZN(_04703_)
);

NAND2_X1 _10347_ (
  .A1(_04702_),
  .A2(_04703_),
  .ZN(_04704_)
);

NAND2_X1 _10348_ (
  .A1(_04704_),
  .A2(_04662_),
  .ZN(_04705_)
);

NAND2_X1 _10349_ (
  .A1(_04675_),
  .A2(\sresult[60][8] ),
  .ZN(_04706_)
);

NAND2_X1 _10350_ (
  .A1(_04705_),
  .A2(_04706_),
  .ZN(_00728_)
);

NAND2_X1 _10351_ (
  .A1(_04670_),
  .A2(\sresult[59][9] ),
  .ZN(_04707_)
);

NAND2_X1 _10352_ (
  .A1(_04659_),
  .A2(din_20[9]),
  .ZN(_04708_)
);

NAND2_X1 _10353_ (
  .A1(_04707_),
  .A2(_04708_),
  .ZN(_04709_)
);

NAND2_X1 _10354_ (
  .A1(_04709_),
  .A2(_04662_),
  .ZN(_04710_)
);

NAND2_X1 _10355_ (
  .A1(_04675_),
  .A2(\sresult[60][9] ),
  .ZN(_04711_)
);

NAND2_X1 _10356_ (
  .A1(_04710_),
  .A2(_04711_),
  .ZN(_00729_)
);

NAND2_X1 _10357_ (
  .A1(_04670_),
  .A2(\sresult[59][10] ),
  .ZN(_04712_)
);

BUF_X4 _10358_ (
  .A(_04279_),
  .Z(_04713_)
);

NAND2_X1 _10359_ (
  .A1(_04713_),
  .A2(din_20[10]),
  .ZN(_04714_)
);

NAND2_X1 _10360_ (
  .A1(_04712_),
  .A2(_04714_),
  .ZN(_04715_)
);

BUF_X1 _10361_ (
  .A(_00911_),
  .Z(_04716_)
);

NAND2_X1 _10362_ (
  .A1(_04715_),
  .A2(_04716_),
  .ZN(_04717_)
);

NAND2_X1 _10363_ (
  .A1(_04675_),
  .A2(\sresult[60][10] ),
  .ZN(_04718_)
);

NAND2_X1 _10364_ (
  .A1(_04717_),
  .A2(_04718_),
  .ZN(_00730_)
);

NAND2_X1 _10365_ (
  .A1(_04670_),
  .A2(\sresult[59][11] ),
  .ZN(_04719_)
);

NAND2_X1 _10366_ (
  .A1(_04713_),
  .A2(din_20[11]),
  .ZN(_04720_)
);

NAND2_X1 _10367_ (
  .A1(_04719_),
  .A2(_04720_),
  .ZN(_04721_)
);

NAND2_X1 _10368_ (
  .A1(_04721_),
  .A2(_04716_),
  .ZN(_04722_)
);

NAND2_X1 _10369_ (
  .A1(_04675_),
  .A2(\sresult[60][11] ),
  .ZN(_04723_)
);

NAND2_X1 _10370_ (
  .A1(_04722_),
  .A2(_04723_),
  .ZN(_00731_)
);

BUF_X4 _10371_ (
  .A(_04235_),
  .Z(_04724_)
);

NAND2_X1 _10372_ (
  .A1(_04724_),
  .A2(\sresult[60][0] ),
  .ZN(_04725_)
);

NAND2_X1 _10373_ (
  .A1(_04713_),
  .A2(din_10[0]),
  .ZN(_04726_)
);

NAND2_X1 _10374_ (
  .A1(_04725_),
  .A2(_04726_),
  .ZN(_04727_)
);

NAND2_X1 _10375_ (
  .A1(_04727_),
  .A2(_04716_),
  .ZN(_04728_)
);

CLKBUF_X2 _10376_ (
  .A(_04296_),
  .Z(_04729_)
);

NAND2_X1 _10377_ (
  .A1(_04729_),
  .A2(\sresult[61][0] ),
  .ZN(_04730_)
);

NAND2_X1 _10378_ (
  .A1(_04728_),
  .A2(_04730_),
  .ZN(_00732_)
);

NAND2_X1 _10379_ (
  .A1(_04724_),
  .A2(\sresult[60][1] ),
  .ZN(_04731_)
);

NAND2_X1 _10380_ (
  .A1(_04713_),
  .A2(din_10[1]),
  .ZN(_04732_)
);

NAND2_X1 _10381_ (
  .A1(_04731_),
  .A2(_04732_),
  .ZN(_04733_)
);

NAND2_X1 _10382_ (
  .A1(_04733_),
  .A2(_04716_),
  .ZN(_04734_)
);

NAND2_X1 _10383_ (
  .A1(_04729_),
  .A2(\sresult[61][1] ),
  .ZN(_04735_)
);

NAND2_X1 _10384_ (
  .A1(_04734_),
  .A2(_04735_),
  .ZN(_00733_)
);

NAND2_X1 _10385_ (
  .A1(_04724_),
  .A2(\sresult[60][2] ),
  .ZN(_04736_)
);

NAND2_X1 _10386_ (
  .A1(_04713_),
  .A2(din_10[2]),
  .ZN(_04737_)
);

NAND2_X1 _10387_ (
  .A1(_04736_),
  .A2(_04737_),
  .ZN(_04738_)
);

NAND2_X1 _10388_ (
  .A1(_04738_),
  .A2(_04716_),
  .ZN(_04739_)
);

NAND2_X1 _10389_ (
  .A1(_04729_),
  .A2(\sresult[61][2] ),
  .ZN(_04740_)
);

NAND2_X1 _10390_ (
  .A1(_04739_),
  .A2(_04740_),
  .ZN(_00734_)
);

NAND2_X1 _10391_ (
  .A1(_04724_),
  .A2(\sresult[60][3] ),
  .ZN(_04741_)
);

NAND2_X1 _10392_ (
  .A1(_04713_),
  .A2(din_10[3]),
  .ZN(_04742_)
);

NAND2_X1 _10393_ (
  .A1(_04741_),
  .A2(_04742_),
  .ZN(_04743_)
);

NAND2_X1 _10394_ (
  .A1(_04743_),
  .A2(_04716_),
  .ZN(_04744_)
);

NAND2_X1 _10395_ (
  .A1(_04729_),
  .A2(\sresult[61][3] ),
  .ZN(_04745_)
);

NAND2_X1 _10396_ (
  .A1(_04744_),
  .A2(_04745_),
  .ZN(_00735_)
);

NAND2_X1 _10397_ (
  .A1(_04724_),
  .A2(\sresult[60][4] ),
  .ZN(_04746_)
);

NAND2_X1 _10398_ (
  .A1(_04713_),
  .A2(din_10[4]),
  .ZN(_04747_)
);

NAND2_X1 _10399_ (
  .A1(_04746_),
  .A2(_04747_),
  .ZN(_04748_)
);

NAND2_X1 _10400_ (
  .A1(_04748_),
  .A2(_04716_),
  .ZN(_04749_)
);

NAND2_X1 _10401_ (
  .A1(_04729_),
  .A2(\sresult[61][4] ),
  .ZN(_04750_)
);

NAND2_X1 _10402_ (
  .A1(_04749_),
  .A2(_04750_),
  .ZN(_00736_)
);

NAND2_X1 _10403_ (
  .A1(_04724_),
  .A2(\sresult[60][5] ),
  .ZN(_04751_)
);

NAND2_X1 _10404_ (
  .A1(_04713_),
  .A2(din_10[5]),
  .ZN(_04752_)
);

NAND2_X1 _10405_ (
  .A1(_04751_),
  .A2(_04752_),
  .ZN(_04753_)
);

NAND2_X1 _10406_ (
  .A1(_04753_),
  .A2(_04716_),
  .ZN(_04754_)
);

NAND2_X1 _10407_ (
  .A1(_04729_),
  .A2(\sresult[61][5] ),
  .ZN(_04755_)
);

NAND2_X1 _10408_ (
  .A1(_04754_),
  .A2(_04755_),
  .ZN(_00737_)
);

NAND2_X1 _10409_ (
  .A1(_04724_),
  .A2(\sresult[60][6] ),
  .ZN(_04756_)
);

NAND2_X1 _10410_ (
  .A1(_04713_),
  .A2(din_10[6]),
  .ZN(_04757_)
);

NAND2_X1 _10411_ (
  .A1(_04756_),
  .A2(_04757_),
  .ZN(_04758_)
);

NAND2_X1 _10412_ (
  .A1(_04758_),
  .A2(_04716_),
  .ZN(_04759_)
);

NAND2_X1 _10413_ (
  .A1(_04729_),
  .A2(\sresult[61][6] ),
  .ZN(_04760_)
);

NAND2_X1 _10414_ (
  .A1(_04759_),
  .A2(_04760_),
  .ZN(_00738_)
);

NAND2_X1 _10415_ (
  .A1(_04724_),
  .A2(\sresult[60][7] ),
  .ZN(_04761_)
);

NAND2_X1 _10416_ (
  .A1(_04713_),
  .A2(din_10[7]),
  .ZN(_04762_)
);

NAND2_X1 _10417_ (
  .A1(_04761_),
  .A2(_04762_),
  .ZN(_04763_)
);

NAND2_X1 _10418_ (
  .A1(_04763_),
  .A2(_04716_),
  .ZN(_04764_)
);

NAND2_X1 _10419_ (
  .A1(_04729_),
  .A2(\sresult[61][7] ),
  .ZN(_04765_)
);

NAND2_X1 _10420_ (
  .A1(_04764_),
  .A2(_04765_),
  .ZN(_00739_)
);

NAND2_X1 _10421_ (
  .A1(_04724_),
  .A2(\sresult[60][8] ),
  .ZN(_04766_)
);

BUF_X4 _10422_ (
  .A(_04279_),
  .Z(_04767_)
);

NAND2_X1 _10423_ (
  .A1(_04767_),
  .A2(din_10[8]),
  .ZN(_04768_)
);

NAND2_X1 _10424_ (
  .A1(_04766_),
  .A2(_04768_),
  .ZN(_04769_)
);

BUF_X1 _10425_ (
  .A(_00911_),
  .Z(_04770_)
);

NAND2_X1 _10426_ (
  .A1(_04769_),
  .A2(_04770_),
  .ZN(_04771_)
);

NAND2_X1 _10427_ (
  .A1(_04729_),
  .A2(\sresult[61][8] ),
  .ZN(_04772_)
);

NAND2_X1 _10428_ (
  .A1(_04771_),
  .A2(_04772_),
  .ZN(_00740_)
);

NAND2_X1 _10429_ (
  .A1(_04724_),
  .A2(\sresult[60][9] ),
  .ZN(_04773_)
);

NAND2_X1 _10430_ (
  .A1(_04767_),
  .A2(din_10[9]),
  .ZN(_04774_)
);

NAND2_X1 _10431_ (
  .A1(_04773_),
  .A2(_04774_),
  .ZN(_04775_)
);

NAND2_X1 _10432_ (
  .A1(_04775_),
  .A2(_04770_),
  .ZN(_04776_)
);

NAND2_X1 _10433_ (
  .A1(_04729_),
  .A2(\sresult[61][9] ),
  .ZN(_04777_)
);

NAND2_X1 _10434_ (
  .A1(_04776_),
  .A2(_04777_),
  .ZN(_00741_)
);

BUF_X2 _10435_ (
  .A(_00799_),
  .Z(_04778_)
);

NAND2_X1 _10436_ (
  .A1(_04778_),
  .A2(\sresult[60][10] ),
  .ZN(_04779_)
);

NAND2_X1 _10437_ (
  .A1(_04767_),
  .A2(din_10[10]),
  .ZN(_04780_)
);

NAND2_X1 _10438_ (
  .A1(_04779_),
  .A2(_04780_),
  .ZN(_04781_)
);

NAND2_X1 _10439_ (
  .A1(_04781_),
  .A2(_04770_),
  .ZN(_04782_)
);

BUF_X2 _10440_ (
  .A(_04296_),
  .Z(_04783_)
);

NAND2_X1 _10441_ (
  .A1(_04783_),
  .A2(\sresult[61][10] ),
  .ZN(_04784_)
);

NAND2_X1 _10442_ (
  .A1(_04782_),
  .A2(_04784_),
  .ZN(_00742_)
);

NAND2_X1 _10443_ (
  .A1(_04778_),
  .A2(\sresult[60][11] ),
  .ZN(_04785_)
);

NAND2_X1 _10444_ (
  .A1(_04767_),
  .A2(din_10[11]),
  .ZN(_04786_)
);

NAND2_X1 _10445_ (
  .A1(_04785_),
  .A2(_04786_),
  .ZN(_04787_)
);

NAND2_X1 _10446_ (
  .A1(_04787_),
  .A2(_04770_),
  .ZN(_04788_)
);

NAND2_X1 _10447_ (
  .A1(_04783_),
  .A2(\sresult[61][11] ),
  .ZN(_04789_)
);

NAND2_X1 _10448_ (
  .A1(_04788_),
  .A2(_04789_),
  .ZN(_00743_)
);

NAND2_X1 _10449_ (
  .A1(_04778_),
  .A2(\sresult[61][0] ),
  .ZN(_04790_)
);

NAND2_X1 _10450_ (
  .A1(_04767_),
  .A2(din_01[0]),
  .ZN(_04791_)
);

NAND2_X1 _10451_ (
  .A1(_04790_),
  .A2(_04791_),
  .ZN(_04792_)
);

NAND2_X1 _10452_ (
  .A1(_04792_),
  .A2(_04770_),
  .ZN(_04793_)
);

NAND2_X1 _10453_ (
  .A1(_04783_),
  .A2(\sresult[62][0] ),
  .ZN(_04794_)
);

NAND2_X1 _10454_ (
  .A1(_04793_),
  .A2(_04794_),
  .ZN(_00744_)
);

NAND2_X1 _10455_ (
  .A1(_04778_),
  .A2(\sresult[61][1] ),
  .ZN(_04795_)
);

NAND2_X1 _10456_ (
  .A1(_04767_),
  .A2(din_01[1]),
  .ZN(_04796_)
);

NAND2_X1 _10457_ (
  .A1(_04795_),
  .A2(_04796_),
  .ZN(_04797_)
);

NAND2_X1 _10458_ (
  .A1(_04797_),
  .A2(_04770_),
  .ZN(_04798_)
);

NAND2_X1 _10459_ (
  .A1(_04783_),
  .A2(\sresult[62][1] ),
  .ZN(_04799_)
);

NAND2_X1 _10460_ (
  .A1(_04798_),
  .A2(_04799_),
  .ZN(_00745_)
);

NAND2_X1 _10461_ (
  .A1(_04778_),
  .A2(\sresult[61][2] ),
  .ZN(_04800_)
);

NAND2_X1 _10462_ (
  .A1(_04767_),
  .A2(din_01[2]),
  .ZN(_04801_)
);

NAND2_X1 _10463_ (
  .A1(_04800_),
  .A2(_04801_),
  .ZN(_04802_)
);

NAND2_X1 _10464_ (
  .A1(_04802_),
  .A2(_04770_),
  .ZN(_04803_)
);

NAND2_X1 _10465_ (
  .A1(_04783_),
  .A2(\sresult[62][2] ),
  .ZN(_04804_)
);

NAND2_X1 _10466_ (
  .A1(_04803_),
  .A2(_04804_),
  .ZN(_00746_)
);

NAND2_X1 _10467_ (
  .A1(_04778_),
  .A2(\sresult[61][3] ),
  .ZN(_04805_)
);

NAND2_X1 _10468_ (
  .A1(_04767_),
  .A2(din_01[3]),
  .ZN(_04806_)
);

NAND2_X1 _10469_ (
  .A1(_04805_),
  .A2(_04806_),
  .ZN(_04807_)
);

NAND2_X1 _10470_ (
  .A1(_04807_),
  .A2(_04770_),
  .ZN(_04808_)
);

NAND2_X1 _10471_ (
  .A1(_04783_),
  .A2(\sresult[62][3] ),
  .ZN(_04809_)
);

NAND2_X1 _10472_ (
  .A1(_04808_),
  .A2(_04809_),
  .ZN(_00747_)
);

NAND2_X1 _10473_ (
  .A1(_04778_),
  .A2(\sresult[61][4] ),
  .ZN(_04810_)
);

NAND2_X1 _10474_ (
  .A1(_04767_),
  .A2(din_01[4]),
  .ZN(_04811_)
);

NAND2_X1 _10475_ (
  .A1(_04810_),
  .A2(_04811_),
  .ZN(_04812_)
);

NAND2_X1 _10476_ (
  .A1(_04812_),
  .A2(_04770_),
  .ZN(_04813_)
);

NAND2_X1 _10477_ (
  .A1(_04783_),
  .A2(\sresult[62][4] ),
  .ZN(_04814_)
);

NAND2_X1 _10478_ (
  .A1(_04813_),
  .A2(_04814_),
  .ZN(_00748_)
);

NAND2_X1 _10479_ (
  .A1(_04778_),
  .A2(\sresult[61][5] ),
  .ZN(_04815_)
);

NAND2_X1 _10480_ (
  .A1(_04767_),
  .A2(din_01[5]),
  .ZN(_04816_)
);

NAND2_X1 _10481_ (
  .A1(_04815_),
  .A2(_04816_),
  .ZN(_04817_)
);

NAND2_X1 _10482_ (
  .A1(_04817_),
  .A2(_04770_),
  .ZN(_04818_)
);

NAND2_X1 _10483_ (
  .A1(_04783_),
  .A2(\sresult[62][5] ),
  .ZN(_04819_)
);

NAND2_X1 _10484_ (
  .A1(_04818_),
  .A2(_04819_),
  .ZN(_00749_)
);

NAND2_X1 _10485_ (
  .A1(_04778_),
  .A2(\sresult[61][6] ),
  .ZN(_04820_)
);

BUF_X2 _10486_ (
  .A(_00770_),
  .Z(_04821_)
);

NAND2_X1 _10487_ (
  .A1(_04821_),
  .A2(din_01[6]),
  .ZN(_04822_)
);

NAND2_X1 _10488_ (
  .A1(_04820_),
  .A2(_04822_),
  .ZN(_04823_)
);

BUF_X1 _10489_ (
  .A(_00911_),
  .Z(_04824_)
);

NAND2_X1 _10490_ (
  .A1(_04823_),
  .A2(_04824_),
  .ZN(_04825_)
);

NAND2_X1 _10491_ (
  .A1(_04783_),
  .A2(\sresult[62][6] ),
  .ZN(_04826_)
);

NAND2_X1 _10492_ (
  .A1(_04825_),
  .A2(_04826_),
  .ZN(_00750_)
);

NAND2_X1 _10493_ (
  .A1(_04778_),
  .A2(\sresult[61][7] ),
  .ZN(_04827_)
);

NAND2_X1 _10494_ (
  .A1(_04821_),
  .A2(din_01[7]),
  .ZN(_04828_)
);

NAND2_X1 _10495_ (
  .A1(_04827_),
  .A2(_04828_),
  .ZN(_04829_)
);

NAND2_X1 _10496_ (
  .A1(_04829_),
  .A2(_04824_),
  .ZN(_04830_)
);

NAND2_X1 _10497_ (
  .A1(_04783_),
  .A2(\sresult[62][7] ),
  .ZN(_04831_)
);

NAND2_X1 _10498_ (
  .A1(_04830_),
  .A2(_04831_),
  .ZN(_00751_)
);

BUF_X2 _10499_ (
  .A(_00799_),
  .Z(_04832_)
);

NAND2_X1 _10500_ (
  .A1(_04832_),
  .A2(\sresult[61][8] ),
  .ZN(_04833_)
);

NAND2_X1 _10501_ (
  .A1(_04821_),
  .A2(din_01[8]),
  .ZN(_04834_)
);

NAND2_X1 _10502_ (
  .A1(_04833_),
  .A2(_04834_),
  .ZN(_04835_)
);

NAND2_X1 _10503_ (
  .A1(_04835_),
  .A2(_04824_),
  .ZN(_04836_)
);

BUF_X1 _10504_ (
  .A(_00810_),
  .Z(_04837_)
);

NAND2_X1 _10505_ (
  .A1(_04837_),
  .A2(\sresult[62][8] ),
  .ZN(_04838_)
);

NAND2_X1 _10506_ (
  .A1(_04836_),
  .A2(_04838_),
  .ZN(_00752_)
);

NAND2_X1 _10507_ (
  .A1(_04832_),
  .A2(\sresult[61][9] ),
  .ZN(_04839_)
);

NAND2_X1 _10508_ (
  .A1(_04821_),
  .A2(din_01[9]),
  .ZN(_04840_)
);

NAND2_X1 _10509_ (
  .A1(_04839_),
  .A2(_04840_),
  .ZN(_04841_)
);

NAND2_X1 _10510_ (
  .A1(_04841_),
  .A2(_04824_),
  .ZN(_04842_)
);

NAND2_X1 _10511_ (
  .A1(_04837_),
  .A2(\sresult[62][9] ),
  .ZN(_04843_)
);

NAND2_X1 _10512_ (
  .A1(_04842_),
  .A2(_04843_),
  .ZN(_00753_)
);

NAND2_X1 _10513_ (
  .A1(_04832_),
  .A2(\sresult[61][10] ),
  .ZN(_04844_)
);

NAND2_X1 _10514_ (
  .A1(_04821_),
  .A2(din_01[10]),
  .ZN(_04845_)
);

NAND2_X1 _10515_ (
  .A1(_04844_),
  .A2(_04845_),
  .ZN(_04846_)
);

NAND2_X1 _10516_ (
  .A1(_04846_),
  .A2(_04824_),
  .ZN(_04847_)
);

NAND2_X1 _10517_ (
  .A1(_04837_),
  .A2(\sresult[62][10] ),
  .ZN(_04848_)
);

NAND2_X1 _10518_ (
  .A1(_04847_),
  .A2(_04848_),
  .ZN(_00754_)
);

NAND2_X1 _10519_ (
  .A1(_04832_),
  .A2(\sresult[61][11] ),
  .ZN(_04849_)
);

NAND2_X1 _10520_ (
  .A1(_04821_),
  .A2(din_01[11]),
  .ZN(_04850_)
);

NAND2_X1 _10521_ (
  .A1(_04849_),
  .A2(_04850_),
  .ZN(_04851_)
);

NAND2_X1 _10522_ (
  .A1(_04851_),
  .A2(_04824_),
  .ZN(_04852_)
);

NAND2_X1 _10523_ (
  .A1(_04837_),
  .A2(\sresult[62][11] ),
  .ZN(_04853_)
);

NAND2_X1 _10524_ (
  .A1(_04852_),
  .A2(_04853_),
  .ZN(_00755_)
);

NAND2_X1 _10525_ (
  .A1(_04832_),
  .A2(\sresult[62][0] ),
  .ZN(_04854_)
);

NAND2_X1 _10526_ (
  .A1(_04821_),
  .A2(din_00[0]),
  .ZN(_04855_)
);

NAND2_X1 _10527_ (
  .A1(_04854_),
  .A2(_04855_),
  .ZN(_04856_)
);

NAND2_X1 _10528_ (
  .A1(_04856_),
  .A2(_04824_),
  .ZN(_04857_)
);

NAND2_X1 _10529_ (
  .A1(_04837_),
  .A2(dout[0]),
  .ZN(_04858_)
);

NAND2_X1 _10530_ (
  .A1(_04857_),
  .A2(_04858_),
  .ZN(_00756_)
);

NAND2_X1 _10531_ (
  .A1(_04832_),
  .A2(\sresult[62][1] ),
  .ZN(_04859_)
);

NAND2_X1 _10532_ (
  .A1(_04821_),
  .A2(din_00[1]),
  .ZN(_04860_)
);

NAND2_X1 _10533_ (
  .A1(_04859_),
  .A2(_04860_),
  .ZN(_04861_)
);

NAND2_X1 _10534_ (
  .A1(_04861_),
  .A2(_04824_),
  .ZN(_04862_)
);

NAND2_X1 _10535_ (
  .A1(_04837_),
  .A2(dout[1]),
  .ZN(_04863_)
);

NAND2_X1 _10536_ (
  .A1(_04862_),
  .A2(_04863_),
  .ZN(_00757_)
);

NAND2_X1 _10537_ (
  .A1(_04832_),
  .A2(\sresult[62][2] ),
  .ZN(_04864_)
);

NAND2_X1 _10538_ (
  .A1(_04821_),
  .A2(din_00[2]),
  .ZN(_04865_)
);

NAND2_X1 _10539_ (
  .A1(_04864_),
  .A2(_04865_),
  .ZN(_04866_)
);

NAND2_X1 _10540_ (
  .A1(_04866_),
  .A2(_04824_),
  .ZN(_04867_)
);

NAND2_X1 _10541_ (
  .A1(_04837_),
  .A2(dout[2]),
  .ZN(_04868_)
);

NAND2_X1 _10542_ (
  .A1(_04867_),
  .A2(_04868_),
  .ZN(_00758_)
);

NAND2_X1 _10543_ (
  .A1(_04832_),
  .A2(\sresult[62][3] ),
  .ZN(_04869_)
);

NAND2_X1 _10544_ (
  .A1(_04821_),
  .A2(din_00[3]),
  .ZN(_04870_)
);

NAND2_X1 _10545_ (
  .A1(_04869_),
  .A2(_04870_),
  .ZN(_04871_)
);

NAND2_X1 _10546_ (
  .A1(_04871_),
  .A2(_04824_),
  .ZN(_04872_)
);

NAND2_X1 _10547_ (
  .A1(_04837_),
  .A2(dout[3]),
  .ZN(_04873_)
);

NAND2_X1 _10548_ (
  .A1(_04872_),
  .A2(_04873_),
  .ZN(_00759_)
);

NAND2_X1 _10549_ (
  .A1(_04832_),
  .A2(\sresult[62][4] ),
  .ZN(_04874_)
);

NAND2_X1 _10550_ (
  .A1(_00803_),
  .A2(din_00[4]),
  .ZN(_04875_)
);

NAND2_X1 _10551_ (
  .A1(_04874_),
  .A2(_04875_),
  .ZN(_04876_)
);

NAND2_X1 _10552_ (
  .A1(_04876_),
  .A2(_00807_),
  .ZN(_04877_)
);

NAND2_X1 _10553_ (
  .A1(_04837_),
  .A2(dout[4]),
  .ZN(_04878_)
);

NAND2_X1 _10554_ (
  .A1(_04877_),
  .A2(_04878_),
  .ZN(_00760_)
);

NAND2_X1 _10555_ (
  .A1(_04832_),
  .A2(\sresult[62][5] ),
  .ZN(_04879_)
);

NAND2_X1 _10556_ (
  .A1(_00803_),
  .A2(din_00[5]),
  .ZN(_04880_)
);

NAND2_X1 _10557_ (
  .A1(_04879_),
  .A2(_04880_),
  .ZN(_04881_)
);

NAND2_X1 _10558_ (
  .A1(_04881_),
  .A2(_00807_),
  .ZN(_04882_)
);

NAND2_X1 _10559_ (
  .A1(_04837_),
  .A2(dout[5]),
  .ZN(_04883_)
);

NAND2_X1 _10560_ (
  .A1(_04882_),
  .A2(_04883_),
  .ZN(_00761_)
);

NAND2_X1 _10561_ (
  .A1(_00814_),
  .A2(\sresult[62][6] ),
  .ZN(_04884_)
);

NAND2_X1 _10562_ (
  .A1(_00803_),
  .A2(din_00[6]),
  .ZN(_04885_)
);

NAND2_X1 _10563_ (
  .A1(_04884_),
  .A2(_04885_),
  .ZN(_04886_)
);

NAND2_X1 _10564_ (
  .A1(_04886_),
  .A2(_00807_),
  .ZN(_04887_)
);

NAND2_X1 _10565_ (
  .A1(_00820_),
  .A2(dout[6]),
  .ZN(_04888_)
);

NAND2_X1 _10566_ (
  .A1(_04887_),
  .A2(_04888_),
  .ZN(_00762_)
);

NAND2_X1 _10567_ (
  .A1(_00814_),
  .A2(\sresult[62][7] ),
  .ZN(_04889_)
);

NAND2_X1 _10568_ (
  .A1(_00803_),
  .A2(din_00[7]),
  .ZN(_04890_)
);

NAND2_X1 _10569_ (
  .A1(_04889_),
  .A2(_04890_),
  .ZN(_04891_)
);

NAND2_X1 _10570_ (
  .A1(_04891_),
  .A2(_00807_),
  .ZN(_04892_)
);

NAND2_X1 _10571_ (
  .A1(_00820_),
  .A2(dout[7]),
  .ZN(_04893_)
);

NAND2_X1 _10572_ (
  .A1(_04892_),
  .A2(_04893_),
  .ZN(_00763_)
);

NAND2_X1 _10573_ (
  .A1(_00814_),
  .A2(\sresult[62][8] ),
  .ZN(_04894_)
);

NAND2_X1 _10574_ (
  .A1(_00804_),
  .A2(din_00[8]),
  .ZN(_04895_)
);

NAND2_X1 _10575_ (
  .A1(_04894_),
  .A2(_04895_),
  .ZN(_04896_)
);

NAND2_X1 _10576_ (
  .A1(_04896_),
  .A2(_00807_),
  .ZN(_04897_)
);

NAND2_X1 _10577_ (
  .A1(_00820_),
  .A2(dout[8]),
  .ZN(_04898_)
);

NAND2_X1 _10578_ (
  .A1(_04897_),
  .A2(_04898_),
  .ZN(_00764_)
);

NAND2_X1 _10579_ (
  .A1(_00814_),
  .A2(\sresult[62][9] ),
  .ZN(_04899_)
);

NAND2_X1 _10580_ (
  .A1(_02813_),
  .A2(din_00[9]),
  .ZN(_04900_)
);

NAND2_X1 _10581_ (
  .A1(_04899_),
  .A2(_04900_),
  .ZN(_04901_)
);

NAND2_X1 _10582_ (
  .A1(_04901_),
  .A2(_00808_),
  .ZN(_04902_)
);

NAND2_X1 _10583_ (
  .A1(_00820_),
  .A2(dout[9]),
  .ZN(_04903_)
);

NAND2_X1 _10584_ (
  .A1(_04902_),
  .A2(_04903_),
  .ZN(_00765_)
);

NAND2_X1 _10585_ (
  .A1(_00814_),
  .A2(\sresult[62][10] ),
  .ZN(_04904_)
);

NAND2_X1 _10586_ (
  .A1(_02813_),
  .A2(din_00[10]),
  .ZN(_04905_)
);

NAND2_X1 _10587_ (
  .A1(_04904_),
  .A2(_04905_),
  .ZN(_04906_)
);

NAND2_X1 _10588_ (
  .A1(_04906_),
  .A2(_02816_),
  .ZN(_04907_)
);

NAND2_X1 _10589_ (
  .A1(_00820_),
  .A2(dout[10]),
  .ZN(_04908_)
);

NAND2_X1 _10590_ (
  .A1(_04907_),
  .A2(_04908_),
  .ZN(_00766_)
);

NAND2_X1 _10591_ (
  .A1(_00814_),
  .A2(\sresult[62][11] ),
  .ZN(_04909_)
);

NAND2_X1 _10592_ (
  .A1(_00804_),
  .A2(din_00[11]),
  .ZN(_04910_)
);

NAND2_X1 _10593_ (
  .A1(_04909_),
  .A2(_04910_),
  .ZN(_04911_)
);

NAND2_X1 _10594_ (
  .A1(_04911_),
  .A2(_02873_),
  .ZN(_04912_)
);

NAND2_X1 _10595_ (
  .A1(_00821_),
  .A2(dout[11]),
  .ZN(_04913_)
);

NAND2_X1 _10596_ (
  .A1(_04912_),
  .A2(_04913_),
  .ZN(_00767_)
);

NAND2_X1 _10597_ (
  .A1(_00807_),
  .A2(dstrb),
  .ZN(_04914_)
);

OAI21_X1 _10598_ (
  .A(_04914_),
  .B1(_00815_),
  .B2(_00808_),
  .ZN(_00768_)
);

DFF_X1 \dout[0]$_DFFE_PP_  (
  .D(_00756_),
  .CK(clk),
  .Q(dout[0]),
  .QN(_04927_)
);

DFF_X1 \dout[10]$_DFFE_PP_  (
  .D(_00766_),
  .CK(clk),
  .Q(dout[10]),
  .QN(_04917_)
);

DFF_X1 \dout[11]$_DFFE_PP_  (
  .D(_00767_),
  .CK(clk),
  .Q(dout[11]),
  .QN(_04916_)
);

DFF_X1 \dout[1]$_DFFE_PP_  (
  .D(_00757_),
  .CK(clk),
  .Q(dout[1]),
  .QN(_04926_)
);

DFF_X1 \dout[2]$_DFFE_PP_  (
  .D(_00758_),
  .CK(clk),
  .Q(dout[2]),
  .QN(_04925_)
);

DFF_X1 \dout[3]$_DFFE_PP_  (
  .D(_00759_),
  .CK(clk),
  .Q(dout[3]),
  .QN(_04924_)
);

DFF_X1 \dout[4]$_DFFE_PP_  (
  .D(_00760_),
  .CK(clk),
  .Q(dout[4]),
  .QN(_04923_)
);

DFF_X1 \dout[5]$_DFFE_PP_  (
  .D(_00761_),
  .CK(clk),
  .Q(dout[5]),
  .QN(_04922_)
);

DFF_X1 \dout[6]$_DFFE_PP_  (
  .D(_00762_),
  .CK(clk),
  .Q(dout[6]),
  .QN(_04921_)
);

DFF_X1 \dout[7]$_DFFE_PP_  (
  .D(_00763_),
  .CK(clk),
  .Q(dout[7]),
  .QN(_04920_)
);

DFF_X1 \dout[8]$_DFFE_PP_  (
  .D(_00764_),
  .CK(clk),
  .Q(dout[8]),
  .QN(_04919_)
);

DFF_X1 \dout[9]$_DFFE_PP_  (
  .D(_00765_),
  .CK(clk),
  .Q(dout[9]),
  .QN(_04918_)
);

DFF_X1 douten$_DFFE_PP_ (
  .D(_00768_),
  .CK(clk),
  .Q(douten),
  .QN(_04915_)
);

DFF_X1 \sresult[0][0]$_DFFE_PP_  (
  .D(_00000_),
  .CK(clk),
  .Q(\sresult[0][0] ),
  .QN(_05683_)
);

DFF_X1 \sresult[0][10]$_DFFE_PP_  (
  .D(_00010_),
  .CK(clk),
  .Q(\sresult[0][10] ),
  .QN(_05673_)
);

DFF_X1 \sresult[0][11]$_DFFE_PP_  (
  .D(_00011_),
  .CK(clk),
  .Q(\sresult[0][11] ),
  .QN(_05672_)
);

DFF_X1 \sresult[0][1]$_DFFE_PP_  (
  .D(_00001_),
  .CK(clk),
  .Q(\sresult[0][1] ),
  .QN(_05682_)
);

DFF_X1 \sresult[0][2]$_DFFE_PP_  (
  .D(_00002_),
  .CK(clk),
  .Q(\sresult[0][2] ),
  .QN(_05681_)
);

DFF_X1 \sresult[0][3]$_DFFE_PP_  (
  .D(_00003_),
  .CK(clk),
  .Q(\sresult[0][3] ),
  .QN(_05680_)
);

DFF_X1 \sresult[0][4]$_DFFE_PP_  (
  .D(_00004_),
  .CK(clk),
  .Q(\sresult[0][4] ),
  .QN(_05679_)
);

DFF_X1 \sresult[0][5]$_DFFE_PP_  (
  .D(_00005_),
  .CK(clk),
  .Q(\sresult[0][5] ),
  .QN(_05678_)
);

DFF_X1 \sresult[0][6]$_DFFE_PP_  (
  .D(_00006_),
  .CK(clk),
  .Q(\sresult[0][6] ),
  .QN(_05677_)
);

DFF_X1 \sresult[0][7]$_DFFE_PP_  (
  .D(_00007_),
  .CK(clk),
  .Q(\sresult[0][7] ),
  .QN(_05676_)
);

DFF_X1 \sresult[0][8]$_DFFE_PP_  (
  .D(_00008_),
  .CK(clk),
  .Q(\sresult[0][8] ),
  .QN(_05675_)
);

DFF_X1 \sresult[0][9]$_DFFE_PP_  (
  .D(_00009_),
  .CK(clk),
  .Q(\sresult[0][9] ),
  .QN(_05674_)
);

DFF_X1 \sresult[10][0]$_DFFE_PP_  (
  .D(_00120_),
  .CK(clk),
  .Q(\sresult[10][0] ),
  .QN(_05563_)
);

DFF_X1 \sresult[10][10]$_DFFE_PP_  (
  .D(_00130_),
  .CK(clk),
  .Q(\sresult[10][10] ),
  .QN(_05553_)
);

DFF_X1 \sresult[10][11]$_DFFE_PP_  (
  .D(_00131_),
  .CK(clk),
  .Q(\sresult[10][11] ),
  .QN(_05552_)
);

DFF_X1 \sresult[10][1]$_DFFE_PP_  (
  .D(_00121_),
  .CK(clk),
  .Q(\sresult[10][1] ),
  .QN(_05562_)
);

DFF_X1 \sresult[10][2]$_DFFE_PP_  (
  .D(_00122_),
  .CK(clk),
  .Q(\sresult[10][2] ),
  .QN(_05561_)
);

DFF_X1 \sresult[10][3]$_DFFE_PP_  (
  .D(_00123_),
  .CK(clk),
  .Q(\sresult[10][3] ),
  .QN(_05560_)
);

DFF_X1 \sresult[10][4]$_DFFE_PP_  (
  .D(_00124_),
  .CK(clk),
  .Q(\sresult[10][4] ),
  .QN(_05559_)
);

DFF_X1 \sresult[10][5]$_DFFE_PP_  (
  .D(_00125_),
  .CK(clk),
  .Q(\sresult[10][5] ),
  .QN(_05558_)
);

DFF_X1 \sresult[10][6]$_DFFE_PP_  (
  .D(_00126_),
  .CK(clk),
  .Q(\sresult[10][6] ),
  .QN(_05557_)
);

DFF_X1 \sresult[10][7]$_DFFE_PP_  (
  .D(_00127_),
  .CK(clk),
  .Q(\sresult[10][7] ),
  .QN(_05556_)
);

DFF_X1 \sresult[10][8]$_DFFE_PP_  (
  .D(_00128_),
  .CK(clk),
  .Q(\sresult[10][8] ),
  .QN(_05555_)
);

DFF_X1 \sresult[10][9]$_DFFE_PP_  (
  .D(_00129_),
  .CK(clk),
  .Q(\sresult[10][9] ),
  .QN(_05554_)
);

DFF_X1 \sresult[11][0]$_DFFE_PP_  (
  .D(_00132_),
  .CK(clk),
  .Q(\sresult[11][0] ),
  .QN(_05551_)
);

DFF_X1 \sresult[11][10]$_DFFE_PP_  (
  .D(_00142_),
  .CK(clk),
  .Q(\sresult[11][10] ),
  .QN(_05541_)
);

DFF_X1 \sresult[11][11]$_DFFE_PP_  (
  .D(_00143_),
  .CK(clk),
  .Q(\sresult[11][11] ),
  .QN(_05540_)
);

DFF_X1 \sresult[11][1]$_DFFE_PP_  (
  .D(_00133_),
  .CK(clk),
  .Q(\sresult[11][1] ),
  .QN(_05550_)
);

DFF_X1 \sresult[11][2]$_DFFE_PP_  (
  .D(_00134_),
  .CK(clk),
  .Q(\sresult[11][2] ),
  .QN(_05549_)
);

DFF_X1 \sresult[11][3]$_DFFE_PP_  (
  .D(_00135_),
  .CK(clk),
  .Q(\sresult[11][3] ),
  .QN(_05548_)
);

DFF_X1 \sresult[11][4]$_DFFE_PP_  (
  .D(_00136_),
  .CK(clk),
  .Q(\sresult[11][4] ),
  .QN(_05547_)
);

DFF_X1 \sresult[11][5]$_DFFE_PP_  (
  .D(_00137_),
  .CK(clk),
  .Q(\sresult[11][5] ),
  .QN(_05546_)
);

DFF_X1 \sresult[11][6]$_DFFE_PP_  (
  .D(_00138_),
  .CK(clk),
  .Q(\sresult[11][6] ),
  .QN(_05545_)
);

DFF_X1 \sresult[11][7]$_DFFE_PP_  (
  .D(_00139_),
  .CK(clk),
  .Q(\sresult[11][7] ),
  .QN(_05544_)
);

DFF_X1 \sresult[11][8]$_DFFE_PP_  (
  .D(_00140_),
  .CK(clk),
  .Q(\sresult[11][8] ),
  .QN(_05543_)
);

DFF_X1 \sresult[11][9]$_DFFE_PP_  (
  .D(_00141_),
  .CK(clk),
  .Q(\sresult[11][9] ),
  .QN(_05542_)
);

DFF_X1 \sresult[12][0]$_DFFE_PP_  (
  .D(_00144_),
  .CK(clk),
  .Q(\sresult[12][0] ),
  .QN(_05539_)
);

DFF_X1 \sresult[12][10]$_DFFE_PP_  (
  .D(_00154_),
  .CK(clk),
  .Q(\sresult[12][10] ),
  .QN(_05529_)
);

DFF_X1 \sresult[12][11]$_DFFE_PP_  (
  .D(_00155_),
  .CK(clk),
  .Q(\sresult[12][11] ),
  .QN(_05528_)
);

DFF_X1 \sresult[12][1]$_DFFE_PP_  (
  .D(_00145_),
  .CK(clk),
  .Q(\sresult[12][1] ),
  .QN(_05538_)
);

DFF_X1 \sresult[12][2]$_DFFE_PP_  (
  .D(_00146_),
  .CK(clk),
  .Q(\sresult[12][2] ),
  .QN(_05537_)
);

DFF_X1 \sresult[12][3]$_DFFE_PP_  (
  .D(_00147_),
  .CK(clk),
  .Q(\sresult[12][3] ),
  .QN(_05536_)
);

DFF_X1 \sresult[12][4]$_DFFE_PP_  (
  .D(_00148_),
  .CK(clk),
  .Q(\sresult[12][4] ),
  .QN(_05535_)
);

DFF_X1 \sresult[12][5]$_DFFE_PP_  (
  .D(_00149_),
  .CK(clk),
  .Q(\sresult[12][5] ),
  .QN(_05534_)
);

DFF_X1 \sresult[12][6]$_DFFE_PP_  (
  .D(_00150_),
  .CK(clk),
  .Q(\sresult[12][6] ),
  .QN(_05533_)
);

DFF_X1 \sresult[12][7]$_DFFE_PP_  (
  .D(_00151_),
  .CK(clk),
  .Q(\sresult[12][7] ),
  .QN(_05532_)
);

DFF_X1 \sresult[12][8]$_DFFE_PP_  (
  .D(_00152_),
  .CK(clk),
  .Q(\sresult[12][8] ),
  .QN(_05531_)
);

DFF_X1 \sresult[12][9]$_DFFE_PP_  (
  .D(_00153_),
  .CK(clk),
  .Q(\sresult[12][9] ),
  .QN(_05530_)
);

DFF_X1 \sresult[13][0]$_DFFE_PP_  (
  .D(_00156_),
  .CK(clk),
  .Q(\sresult[13][0] ),
  .QN(_05527_)
);

DFF_X1 \sresult[13][10]$_DFFE_PP_  (
  .D(_00166_),
  .CK(clk),
  .Q(\sresult[13][10] ),
  .QN(_05517_)
);

DFF_X1 \sresult[13][11]$_DFFE_PP_  (
  .D(_00167_),
  .CK(clk),
  .Q(\sresult[13][11] ),
  .QN(_05516_)
);

DFF_X1 \sresult[13][1]$_DFFE_PP_  (
  .D(_00157_),
  .CK(clk),
  .Q(\sresult[13][1] ),
  .QN(_05526_)
);

DFF_X1 \sresult[13][2]$_DFFE_PP_  (
  .D(_00158_),
  .CK(clk),
  .Q(\sresult[13][2] ),
  .QN(_05525_)
);

DFF_X1 \sresult[13][3]$_DFFE_PP_  (
  .D(_00159_),
  .CK(clk),
  .Q(\sresult[13][3] ),
  .QN(_05524_)
);

DFF_X1 \sresult[13][4]$_DFFE_PP_  (
  .D(_00160_),
  .CK(clk),
  .Q(\sresult[13][4] ),
  .QN(_05523_)
);

DFF_X1 \sresult[13][5]$_DFFE_PP_  (
  .D(_00161_),
  .CK(clk),
  .Q(\sresult[13][5] ),
  .QN(_05522_)
);

DFF_X1 \sresult[13][6]$_DFFE_PP_  (
  .D(_00162_),
  .CK(clk),
  .Q(\sresult[13][6] ),
  .QN(_05521_)
);

DFF_X1 \sresult[13][7]$_DFFE_PP_  (
  .D(_00163_),
  .CK(clk),
  .Q(\sresult[13][7] ),
  .QN(_05520_)
);

DFF_X1 \sresult[13][8]$_DFFE_PP_  (
  .D(_00164_),
  .CK(clk),
  .Q(\sresult[13][8] ),
  .QN(_05519_)
);

DFF_X1 \sresult[13][9]$_DFFE_PP_  (
  .D(_00165_),
  .CK(clk),
  .Q(\sresult[13][9] ),
  .QN(_05518_)
);

DFF_X1 \sresult[14][0]$_DFFE_PP_  (
  .D(_00168_),
  .CK(clk),
  .Q(\sresult[14][0] ),
  .QN(_05515_)
);

DFF_X1 \sresult[14][10]$_DFFE_PP_  (
  .D(_00178_),
  .CK(clk),
  .Q(\sresult[14][10] ),
  .QN(_05505_)
);

DFF_X1 \sresult[14][11]$_DFFE_PP_  (
  .D(_00179_),
  .CK(clk),
  .Q(\sresult[14][11] ),
  .QN(_05504_)
);

DFF_X1 \sresult[14][1]$_DFFE_PP_  (
  .D(_00169_),
  .CK(clk),
  .Q(\sresult[14][1] ),
  .QN(_05514_)
);

DFF_X1 \sresult[14][2]$_DFFE_PP_  (
  .D(_00170_),
  .CK(clk),
  .Q(\sresult[14][2] ),
  .QN(_05513_)
);

DFF_X1 \sresult[14][3]$_DFFE_PP_  (
  .D(_00171_),
  .CK(clk),
  .Q(\sresult[14][3] ),
  .QN(_05512_)
);

DFF_X1 \sresult[14][4]$_DFFE_PP_  (
  .D(_00172_),
  .CK(clk),
  .Q(\sresult[14][4] ),
  .QN(_05511_)
);

DFF_X1 \sresult[14][5]$_DFFE_PP_  (
  .D(_00173_),
  .CK(clk),
  .Q(\sresult[14][5] ),
  .QN(_05510_)
);

DFF_X1 \sresult[14][6]$_DFFE_PP_  (
  .D(_00174_),
  .CK(clk),
  .Q(\sresult[14][6] ),
  .QN(_05509_)
);

DFF_X1 \sresult[14][7]$_DFFE_PP_  (
  .D(_00175_),
  .CK(clk),
  .Q(\sresult[14][7] ),
  .QN(_05508_)
);

DFF_X1 \sresult[14][8]$_DFFE_PP_  (
  .D(_00176_),
  .CK(clk),
  .Q(\sresult[14][8] ),
  .QN(_05507_)
);

DFF_X1 \sresult[14][9]$_DFFE_PP_  (
  .D(_00177_),
  .CK(clk),
  .Q(\sresult[14][9] ),
  .QN(_05506_)
);

DFF_X1 \sresult[15][0]$_DFFE_PP_  (
  .D(_00180_),
  .CK(clk),
  .Q(\sresult[15][0] ),
  .QN(_05503_)
);

DFF_X1 \sresult[15][10]$_DFFE_PP_  (
  .D(_00190_),
  .CK(clk),
  .Q(\sresult[15][10] ),
  .QN(_05493_)
);

DFF_X1 \sresult[15][11]$_DFFE_PP_  (
  .D(_00191_),
  .CK(clk),
  .Q(\sresult[15][11] ),
  .QN(_05492_)
);

DFF_X1 \sresult[15][1]$_DFFE_PP_  (
  .D(_00181_),
  .CK(clk),
  .Q(\sresult[15][1] ),
  .QN(_05502_)
);

DFF_X1 \sresult[15][2]$_DFFE_PP_  (
  .D(_00182_),
  .CK(clk),
  .Q(\sresult[15][2] ),
  .QN(_05501_)
);

DFF_X1 \sresult[15][3]$_DFFE_PP_  (
  .D(_00183_),
  .CK(clk),
  .Q(\sresult[15][3] ),
  .QN(_05500_)
);

DFF_X1 \sresult[15][4]$_DFFE_PP_  (
  .D(_00184_),
  .CK(clk),
  .Q(\sresult[15][4] ),
  .QN(_05499_)
);

DFF_X1 \sresult[15][5]$_DFFE_PP_  (
  .D(_00185_),
  .CK(clk),
  .Q(\sresult[15][5] ),
  .QN(_05498_)
);

DFF_X1 \sresult[15][6]$_DFFE_PP_  (
  .D(_00186_),
  .CK(clk),
  .Q(\sresult[15][6] ),
  .QN(_05497_)
);

DFF_X1 \sresult[15][7]$_DFFE_PP_  (
  .D(_00187_),
  .CK(clk),
  .Q(\sresult[15][7] ),
  .QN(_05496_)
);

DFF_X1 \sresult[15][8]$_DFFE_PP_  (
  .D(_00188_),
  .CK(clk),
  .Q(\sresult[15][8] ),
  .QN(_05495_)
);

DFF_X1 \sresult[15][9]$_DFFE_PP_  (
  .D(_00189_),
  .CK(clk),
  .Q(\sresult[15][9] ),
  .QN(_05494_)
);

DFF_X1 \sresult[16][0]$_DFFE_PP_  (
  .D(_00192_),
  .CK(clk),
  .Q(\sresult[16][0] ),
  .QN(_05491_)
);

DFF_X1 \sresult[16][10]$_DFFE_PP_  (
  .D(_00202_),
  .CK(clk),
  .Q(\sresult[16][10] ),
  .QN(_05481_)
);

DFF_X1 \sresult[16][11]$_DFFE_PP_  (
  .D(_00203_),
  .CK(clk),
  .Q(\sresult[16][11] ),
  .QN(_05480_)
);

DFF_X1 \sresult[16][1]$_DFFE_PP_  (
  .D(_00193_),
  .CK(clk),
  .Q(\sresult[16][1] ),
  .QN(_05490_)
);

DFF_X1 \sresult[16][2]$_DFFE_PP_  (
  .D(_00194_),
  .CK(clk),
  .Q(\sresult[16][2] ),
  .QN(_05489_)
);

DFF_X1 \sresult[16][3]$_DFFE_PP_  (
  .D(_00195_),
  .CK(clk),
  .Q(\sresult[16][3] ),
  .QN(_05488_)
);

DFF_X1 \sresult[16][4]$_DFFE_PP_  (
  .D(_00196_),
  .CK(clk),
  .Q(\sresult[16][4] ),
  .QN(_05487_)
);

DFF_X1 \sresult[16][5]$_DFFE_PP_  (
  .D(_00197_),
  .CK(clk),
  .Q(\sresult[16][5] ),
  .QN(_05486_)
);

DFF_X1 \sresult[16][6]$_DFFE_PP_  (
  .D(_00198_),
  .CK(clk),
  .Q(\sresult[16][6] ),
  .QN(_05485_)
);

DFF_X1 \sresult[16][7]$_DFFE_PP_  (
  .D(_00199_),
  .CK(clk),
  .Q(\sresult[16][7] ),
  .QN(_05484_)
);

DFF_X1 \sresult[16][8]$_DFFE_PP_  (
  .D(_00200_),
  .CK(clk),
  .Q(\sresult[16][8] ),
  .QN(_05483_)
);

DFF_X1 \sresult[16][9]$_DFFE_PP_  (
  .D(_00201_),
  .CK(clk),
  .Q(\sresult[16][9] ),
  .QN(_05482_)
);

DFF_X1 \sresult[17][0]$_DFFE_PP_  (
  .D(_00204_),
  .CK(clk),
  .Q(\sresult[17][0] ),
  .QN(_05479_)
);

DFF_X1 \sresult[17][10]$_DFFE_PP_  (
  .D(_00214_),
  .CK(clk),
  .Q(\sresult[17][10] ),
  .QN(_05469_)
);

DFF_X1 \sresult[17][11]$_DFFE_PP_  (
  .D(_00215_),
  .CK(clk),
  .Q(\sresult[17][11] ),
  .QN(_05468_)
);

DFF_X1 \sresult[17][1]$_DFFE_PP_  (
  .D(_00205_),
  .CK(clk),
  .Q(\sresult[17][1] ),
  .QN(_05478_)
);

DFF_X1 \sresult[17][2]$_DFFE_PP_  (
  .D(_00206_),
  .CK(clk),
  .Q(\sresult[17][2] ),
  .QN(_05477_)
);

DFF_X1 \sresult[17][3]$_DFFE_PP_  (
  .D(_00207_),
  .CK(clk),
  .Q(\sresult[17][3] ),
  .QN(_05476_)
);

DFF_X1 \sresult[17][4]$_DFFE_PP_  (
  .D(_00208_),
  .CK(clk),
  .Q(\sresult[17][4] ),
  .QN(_05475_)
);

DFF_X1 \sresult[17][5]$_DFFE_PP_  (
  .D(_00209_),
  .CK(clk),
  .Q(\sresult[17][5] ),
  .QN(_05474_)
);

DFF_X1 \sresult[17][6]$_DFFE_PP_  (
  .D(_00210_),
  .CK(clk),
  .Q(\sresult[17][6] ),
  .QN(_05473_)
);

DFF_X1 \sresult[17][7]$_DFFE_PP_  (
  .D(_00211_),
  .CK(clk),
  .Q(\sresult[17][7] ),
  .QN(_05472_)
);

DFF_X1 \sresult[17][8]$_DFFE_PP_  (
  .D(_00212_),
  .CK(clk),
  .Q(\sresult[17][8] ),
  .QN(_05471_)
);

DFF_X1 \sresult[17][9]$_DFFE_PP_  (
  .D(_00213_),
  .CK(clk),
  .Q(\sresult[17][9] ),
  .QN(_05470_)
);

DFF_X1 \sresult[18][0]$_DFFE_PP_  (
  .D(_00216_),
  .CK(clk),
  .Q(\sresult[18][0] ),
  .QN(_05467_)
);

DFF_X1 \sresult[18][10]$_DFFE_PP_  (
  .D(_00226_),
  .CK(clk),
  .Q(\sresult[18][10] ),
  .QN(_05457_)
);

DFF_X1 \sresult[18][11]$_DFFE_PP_  (
  .D(_00227_),
  .CK(clk),
  .Q(\sresult[18][11] ),
  .QN(_05456_)
);

DFF_X1 \sresult[18][1]$_DFFE_PP_  (
  .D(_00217_),
  .CK(clk),
  .Q(\sresult[18][1] ),
  .QN(_05466_)
);

DFF_X1 \sresult[18][2]$_DFFE_PP_  (
  .D(_00218_),
  .CK(clk),
  .Q(\sresult[18][2] ),
  .QN(_05465_)
);

DFF_X1 \sresult[18][3]$_DFFE_PP_  (
  .D(_00219_),
  .CK(clk),
  .Q(\sresult[18][3] ),
  .QN(_05464_)
);

DFF_X1 \sresult[18][4]$_DFFE_PP_  (
  .D(_00220_),
  .CK(clk),
  .Q(\sresult[18][4] ),
  .QN(_05463_)
);

DFF_X1 \sresult[18][5]$_DFFE_PP_  (
  .D(_00221_),
  .CK(clk),
  .Q(\sresult[18][5] ),
  .QN(_05462_)
);

DFF_X1 \sresult[18][6]$_DFFE_PP_  (
  .D(_00222_),
  .CK(clk),
  .Q(\sresult[18][6] ),
  .QN(_05461_)
);

DFF_X1 \sresult[18][7]$_DFFE_PP_  (
  .D(_00223_),
  .CK(clk),
  .Q(\sresult[18][7] ),
  .QN(_05460_)
);

DFF_X1 \sresult[18][8]$_DFFE_PP_  (
  .D(_00224_),
  .CK(clk),
  .Q(\sresult[18][8] ),
  .QN(_05459_)
);

DFF_X1 \sresult[18][9]$_DFFE_PP_  (
  .D(_00225_),
  .CK(clk),
  .Q(\sresult[18][9] ),
  .QN(_05458_)
);

DFF_X1 \sresult[19][0]$_DFFE_PP_  (
  .D(_00228_),
  .CK(clk),
  .Q(\sresult[19][0] ),
  .QN(_05455_)
);

DFF_X1 \sresult[19][10]$_DFFE_PP_  (
  .D(_00238_),
  .CK(clk),
  .Q(\sresult[19][10] ),
  .QN(_05445_)
);

DFF_X1 \sresult[19][11]$_DFFE_PP_  (
  .D(_00239_),
  .CK(clk),
  .Q(\sresult[19][11] ),
  .QN(_05444_)
);

DFF_X1 \sresult[19][1]$_DFFE_PP_  (
  .D(_00229_),
  .CK(clk),
  .Q(\sresult[19][1] ),
  .QN(_05454_)
);

DFF_X1 \sresult[19][2]$_DFFE_PP_  (
  .D(_00230_),
  .CK(clk),
  .Q(\sresult[19][2] ),
  .QN(_05453_)
);

DFF_X1 \sresult[19][3]$_DFFE_PP_  (
  .D(_00231_),
  .CK(clk),
  .Q(\sresult[19][3] ),
  .QN(_05452_)
);

DFF_X1 \sresult[19][4]$_DFFE_PP_  (
  .D(_00232_),
  .CK(clk),
  .Q(\sresult[19][4] ),
  .QN(_05451_)
);

DFF_X1 \sresult[19][5]$_DFFE_PP_  (
  .D(_00233_),
  .CK(clk),
  .Q(\sresult[19][5] ),
  .QN(_05450_)
);

DFF_X1 \sresult[19][6]$_DFFE_PP_  (
  .D(_00234_),
  .CK(clk),
  .Q(\sresult[19][6] ),
  .QN(_05449_)
);

DFF_X1 \sresult[19][7]$_DFFE_PP_  (
  .D(_00235_),
  .CK(clk),
  .Q(\sresult[19][7] ),
  .QN(_05448_)
);

DFF_X1 \sresult[19][8]$_DFFE_PP_  (
  .D(_00236_),
  .CK(clk),
  .Q(\sresult[19][8] ),
  .QN(_05447_)
);

DFF_X1 \sresult[19][9]$_DFFE_PP_  (
  .D(_00237_),
  .CK(clk),
  .Q(\sresult[19][9] ),
  .QN(_05446_)
);

DFF_X1 \sresult[1][0]$_DFFE_PP_  (
  .D(_00012_),
  .CK(clk),
  .Q(\sresult[1][0] ),
  .QN(_05671_)
);

DFF_X1 \sresult[1][10]$_DFFE_PP_  (
  .D(_00022_),
  .CK(clk),
  .Q(\sresult[1][10] ),
  .QN(_05661_)
);

DFF_X1 \sresult[1][11]$_DFFE_PP_  (
  .D(_00023_),
  .CK(clk),
  .Q(\sresult[1][11] ),
  .QN(_05660_)
);

DFF_X1 \sresult[1][1]$_DFFE_PP_  (
  .D(_00013_),
  .CK(clk),
  .Q(\sresult[1][1] ),
  .QN(_05670_)
);

DFF_X1 \sresult[1][2]$_DFFE_PP_  (
  .D(_00014_),
  .CK(clk),
  .Q(\sresult[1][2] ),
  .QN(_05669_)
);

DFF_X1 \sresult[1][3]$_DFFE_PP_  (
  .D(_00015_),
  .CK(clk),
  .Q(\sresult[1][3] ),
  .QN(_05668_)
);

DFF_X1 \sresult[1][4]$_DFFE_PP_  (
  .D(_00016_),
  .CK(clk),
  .Q(\sresult[1][4] ),
  .QN(_05667_)
);

DFF_X1 \sresult[1][5]$_DFFE_PP_  (
  .D(_00017_),
  .CK(clk),
  .Q(\sresult[1][5] ),
  .QN(_05666_)
);

DFF_X1 \sresult[1][6]$_DFFE_PP_  (
  .D(_00018_),
  .CK(clk),
  .Q(\sresult[1][6] ),
  .QN(_05665_)
);

DFF_X1 \sresult[1][7]$_DFFE_PP_  (
  .D(_00019_),
  .CK(clk),
  .Q(\sresult[1][7] ),
  .QN(_05664_)
);

DFF_X1 \sresult[1][8]$_DFFE_PP_  (
  .D(_00020_),
  .CK(clk),
  .Q(\sresult[1][8] ),
  .QN(_05663_)
);

DFF_X1 \sresult[1][9]$_DFFE_PP_  (
  .D(_00021_),
  .CK(clk),
  .Q(\sresult[1][9] ),
  .QN(_05662_)
);

DFF_X1 \sresult[20][0]$_DFFE_PP_  (
  .D(_00240_),
  .CK(clk),
  .Q(\sresult[20][0] ),
  .QN(_05443_)
);

DFF_X1 \sresult[20][10]$_DFFE_PP_  (
  .D(_00250_),
  .CK(clk),
  .Q(\sresult[20][10] ),
  .QN(_05433_)
);

DFF_X1 \sresult[20][11]$_DFFE_PP_  (
  .D(_00251_),
  .CK(clk),
  .Q(\sresult[20][11] ),
  .QN(_05432_)
);

DFF_X1 \sresult[20][1]$_DFFE_PP_  (
  .D(_00241_),
  .CK(clk),
  .Q(\sresult[20][1] ),
  .QN(_05442_)
);

DFF_X1 \sresult[20][2]$_DFFE_PP_  (
  .D(_00242_),
  .CK(clk),
  .Q(\sresult[20][2] ),
  .QN(_05441_)
);

DFF_X1 \sresult[20][3]$_DFFE_PP_  (
  .D(_00243_),
  .CK(clk),
  .Q(\sresult[20][3] ),
  .QN(_05440_)
);

DFF_X1 \sresult[20][4]$_DFFE_PP_  (
  .D(_00244_),
  .CK(clk),
  .Q(\sresult[20][4] ),
  .QN(_05439_)
);

DFF_X1 \sresult[20][5]$_DFFE_PP_  (
  .D(_00245_),
  .CK(clk),
  .Q(\sresult[20][5] ),
  .QN(_05438_)
);

DFF_X1 \sresult[20][6]$_DFFE_PP_  (
  .D(_00246_),
  .CK(clk),
  .Q(\sresult[20][6] ),
  .QN(_05437_)
);

DFF_X1 \sresult[20][7]$_DFFE_PP_  (
  .D(_00247_),
  .CK(clk),
  .Q(\sresult[20][7] ),
  .QN(_05436_)
);

DFF_X1 \sresult[20][8]$_DFFE_PP_  (
  .D(_00248_),
  .CK(clk),
  .Q(\sresult[20][8] ),
  .QN(_05435_)
);

DFF_X1 \sresult[20][9]$_DFFE_PP_  (
  .D(_00249_),
  .CK(clk),
  .Q(\sresult[20][9] ),
  .QN(_05434_)
);

DFF_X1 \sresult[21][0]$_DFFE_PP_  (
  .D(_00252_),
  .CK(clk),
  .Q(\sresult[21][0] ),
  .QN(_05431_)
);

DFF_X1 \sresult[21][10]$_DFFE_PP_  (
  .D(_00262_),
  .CK(clk),
  .Q(\sresult[21][10] ),
  .QN(_05421_)
);

DFF_X1 \sresult[21][11]$_DFFE_PP_  (
  .D(_00263_),
  .CK(clk),
  .Q(\sresult[21][11] ),
  .QN(_05420_)
);

DFF_X1 \sresult[21][1]$_DFFE_PP_  (
  .D(_00253_),
  .CK(clk),
  .Q(\sresult[21][1] ),
  .QN(_05430_)
);

DFF_X1 \sresult[21][2]$_DFFE_PP_  (
  .D(_00254_),
  .CK(clk),
  .Q(\sresult[21][2] ),
  .QN(_05429_)
);

DFF_X1 \sresult[21][3]$_DFFE_PP_  (
  .D(_00255_),
  .CK(clk),
  .Q(\sresult[21][3] ),
  .QN(_05428_)
);

DFF_X1 \sresult[21][4]$_DFFE_PP_  (
  .D(_00256_),
  .CK(clk),
  .Q(\sresult[21][4] ),
  .QN(_05427_)
);

DFF_X1 \sresult[21][5]$_DFFE_PP_  (
  .D(_00257_),
  .CK(clk),
  .Q(\sresult[21][5] ),
  .QN(_05426_)
);

DFF_X1 \sresult[21][6]$_DFFE_PP_  (
  .D(_00258_),
  .CK(clk),
  .Q(\sresult[21][6] ),
  .QN(_05425_)
);

DFF_X1 \sresult[21][7]$_DFFE_PP_  (
  .D(_00259_),
  .CK(clk),
  .Q(\sresult[21][7] ),
  .QN(_05424_)
);

DFF_X1 \sresult[21][8]$_DFFE_PP_  (
  .D(_00260_),
  .CK(clk),
  .Q(\sresult[21][8] ),
  .QN(_05423_)
);

DFF_X1 \sresult[21][9]$_DFFE_PP_  (
  .D(_00261_),
  .CK(clk),
  .Q(\sresult[21][9] ),
  .QN(_05422_)
);

DFF_X1 \sresult[22][0]$_DFFE_PP_  (
  .D(_00264_),
  .CK(clk),
  .Q(\sresult[22][0] ),
  .QN(_05419_)
);

DFF_X1 \sresult[22][10]$_DFFE_PP_  (
  .D(_00274_),
  .CK(clk),
  .Q(\sresult[22][10] ),
  .QN(_05409_)
);

DFF_X1 \sresult[22][11]$_DFFE_PP_  (
  .D(_00275_),
  .CK(clk),
  .Q(\sresult[22][11] ),
  .QN(_05408_)
);

DFF_X1 \sresult[22][1]$_DFFE_PP_  (
  .D(_00265_),
  .CK(clk),
  .Q(\sresult[22][1] ),
  .QN(_05418_)
);

DFF_X1 \sresult[22][2]$_DFFE_PP_  (
  .D(_00266_),
  .CK(clk),
  .Q(\sresult[22][2] ),
  .QN(_05417_)
);

DFF_X1 \sresult[22][3]$_DFFE_PP_  (
  .D(_00267_),
  .CK(clk),
  .Q(\sresult[22][3] ),
  .QN(_05416_)
);

DFF_X1 \sresult[22][4]$_DFFE_PP_  (
  .D(_00268_),
  .CK(clk),
  .Q(\sresult[22][4] ),
  .QN(_05415_)
);

DFF_X1 \sresult[22][5]$_DFFE_PP_  (
  .D(_00269_),
  .CK(clk),
  .Q(\sresult[22][5] ),
  .QN(_05414_)
);

DFF_X1 \sresult[22][6]$_DFFE_PP_  (
  .D(_00270_),
  .CK(clk),
  .Q(\sresult[22][6] ),
  .QN(_05413_)
);

DFF_X1 \sresult[22][7]$_DFFE_PP_  (
  .D(_00271_),
  .CK(clk),
  .Q(\sresult[22][7] ),
  .QN(_05412_)
);

DFF_X1 \sresult[22][8]$_DFFE_PP_  (
  .D(_00272_),
  .CK(clk),
  .Q(\sresult[22][8] ),
  .QN(_05411_)
);

DFF_X1 \sresult[22][9]$_DFFE_PP_  (
  .D(_00273_),
  .CK(clk),
  .Q(\sresult[22][9] ),
  .QN(_05410_)
);

DFF_X1 \sresult[23][0]$_DFFE_PP_  (
  .D(_00276_),
  .CK(clk),
  .Q(\sresult[23][0] ),
  .QN(_05407_)
);

DFF_X1 \sresult[23][10]$_DFFE_PP_  (
  .D(_00286_),
  .CK(clk),
  .Q(\sresult[23][10] ),
  .QN(_05397_)
);

DFF_X1 \sresult[23][11]$_DFFE_PP_  (
  .D(_00287_),
  .CK(clk),
  .Q(\sresult[23][11] ),
  .QN(_05396_)
);

DFF_X1 \sresult[23][1]$_DFFE_PP_  (
  .D(_00277_),
  .CK(clk),
  .Q(\sresult[23][1] ),
  .QN(_05406_)
);

DFF_X1 \sresult[23][2]$_DFFE_PP_  (
  .D(_00278_),
  .CK(clk),
  .Q(\sresult[23][2] ),
  .QN(_05405_)
);

DFF_X1 \sresult[23][3]$_DFFE_PP_  (
  .D(_00279_),
  .CK(clk),
  .Q(\sresult[23][3] ),
  .QN(_05404_)
);

DFF_X1 \sresult[23][4]$_DFFE_PP_  (
  .D(_00280_),
  .CK(clk),
  .Q(\sresult[23][4] ),
  .QN(_05403_)
);

DFF_X1 \sresult[23][5]$_DFFE_PP_  (
  .D(_00281_),
  .CK(clk),
  .Q(\sresult[23][5] ),
  .QN(_05402_)
);

DFF_X1 \sresult[23][6]$_DFFE_PP_  (
  .D(_00282_),
  .CK(clk),
  .Q(\sresult[23][6] ),
  .QN(_05401_)
);

DFF_X1 \sresult[23][7]$_DFFE_PP_  (
  .D(_00283_),
  .CK(clk),
  .Q(\sresult[23][7] ),
  .QN(_05400_)
);

DFF_X1 \sresult[23][8]$_DFFE_PP_  (
  .D(_00284_),
  .CK(clk),
  .Q(\sresult[23][8] ),
  .QN(_05399_)
);

DFF_X1 \sresult[23][9]$_DFFE_PP_  (
  .D(_00285_),
  .CK(clk),
  .Q(\sresult[23][9] ),
  .QN(_05398_)
);

DFF_X1 \sresult[24][0]$_DFFE_PP_  (
  .D(_00288_),
  .CK(clk),
  .Q(\sresult[24][0] ),
  .QN(_05395_)
);

DFF_X1 \sresult[24][10]$_DFFE_PP_  (
  .D(_00298_),
  .CK(clk),
  .Q(\sresult[24][10] ),
  .QN(_05385_)
);

DFF_X1 \sresult[24][11]$_DFFE_PP_  (
  .D(_00299_),
  .CK(clk),
  .Q(\sresult[24][11] ),
  .QN(_05384_)
);

DFF_X1 \sresult[24][1]$_DFFE_PP_  (
  .D(_00289_),
  .CK(clk),
  .Q(\sresult[24][1] ),
  .QN(_05394_)
);

DFF_X1 \sresult[24][2]$_DFFE_PP_  (
  .D(_00290_),
  .CK(clk),
  .Q(\sresult[24][2] ),
  .QN(_05393_)
);

DFF_X1 \sresult[24][3]$_DFFE_PP_  (
  .D(_00291_),
  .CK(clk),
  .Q(\sresult[24][3] ),
  .QN(_05392_)
);

DFF_X1 \sresult[24][4]$_DFFE_PP_  (
  .D(_00292_),
  .CK(clk),
  .Q(\sresult[24][4] ),
  .QN(_05391_)
);

DFF_X1 \sresult[24][5]$_DFFE_PP_  (
  .D(_00293_),
  .CK(clk),
  .Q(\sresult[24][5] ),
  .QN(_05390_)
);

DFF_X1 \sresult[24][6]$_DFFE_PP_  (
  .D(_00294_),
  .CK(clk),
  .Q(\sresult[24][6] ),
  .QN(_05389_)
);

DFF_X1 \sresult[24][7]$_DFFE_PP_  (
  .D(_00295_),
  .CK(clk),
  .Q(\sresult[24][7] ),
  .QN(_05388_)
);

DFF_X1 \sresult[24][8]$_DFFE_PP_  (
  .D(_00296_),
  .CK(clk),
  .Q(\sresult[24][8] ),
  .QN(_05387_)
);

DFF_X1 \sresult[24][9]$_DFFE_PP_  (
  .D(_00297_),
  .CK(clk),
  .Q(\sresult[24][9] ),
  .QN(_05386_)
);

DFF_X1 \sresult[25][0]$_DFFE_PP_  (
  .D(_00300_),
  .CK(clk),
  .Q(\sresult[25][0] ),
  .QN(_05383_)
);

DFF_X1 \sresult[25][10]$_DFFE_PP_  (
  .D(_00310_),
  .CK(clk),
  .Q(\sresult[25][10] ),
  .QN(_05373_)
);

DFF_X1 \sresult[25][11]$_DFFE_PP_  (
  .D(_00311_),
  .CK(clk),
  .Q(\sresult[25][11] ),
  .QN(_05372_)
);

DFF_X1 \sresult[25][1]$_DFFE_PP_  (
  .D(_00301_),
  .CK(clk),
  .Q(\sresult[25][1] ),
  .QN(_05382_)
);

DFF_X1 \sresult[25][2]$_DFFE_PP_  (
  .D(_00302_),
  .CK(clk),
  .Q(\sresult[25][2] ),
  .QN(_05381_)
);

DFF_X1 \sresult[25][3]$_DFFE_PP_  (
  .D(_00303_),
  .CK(clk),
  .Q(\sresult[25][3] ),
  .QN(_05380_)
);

DFF_X1 \sresult[25][4]$_DFFE_PP_  (
  .D(_00304_),
  .CK(clk),
  .Q(\sresult[25][4] ),
  .QN(_05379_)
);

DFF_X1 \sresult[25][5]$_DFFE_PP_  (
  .D(_00305_),
  .CK(clk),
  .Q(\sresult[25][5] ),
  .QN(_05378_)
);

DFF_X1 \sresult[25][6]$_DFFE_PP_  (
  .D(_00306_),
  .CK(clk),
  .Q(\sresult[25][6] ),
  .QN(_05377_)
);

DFF_X1 \sresult[25][7]$_DFFE_PP_  (
  .D(_00307_),
  .CK(clk),
  .Q(\sresult[25][7] ),
  .QN(_05376_)
);

DFF_X1 \sresult[25][8]$_DFFE_PP_  (
  .D(_00308_),
  .CK(clk),
  .Q(\sresult[25][8] ),
  .QN(_05375_)
);

DFF_X1 \sresult[25][9]$_DFFE_PP_  (
  .D(_00309_),
  .CK(clk),
  .Q(\sresult[25][9] ),
  .QN(_05374_)
);

DFF_X1 \sresult[26][0]$_DFFE_PP_  (
  .D(_00312_),
  .CK(clk),
  .Q(\sresult[26][0] ),
  .QN(_05371_)
);

DFF_X1 \sresult[26][10]$_DFFE_PP_  (
  .D(_00322_),
  .CK(clk),
  .Q(\sresult[26][10] ),
  .QN(_05361_)
);

DFF_X1 \sresult[26][11]$_DFFE_PP_  (
  .D(_00323_),
  .CK(clk),
  .Q(\sresult[26][11] ),
  .QN(_05360_)
);

DFF_X1 \sresult[26][1]$_DFFE_PP_  (
  .D(_00313_),
  .CK(clk),
  .Q(\sresult[26][1] ),
  .QN(_05370_)
);

DFF_X1 \sresult[26][2]$_DFFE_PP_  (
  .D(_00314_),
  .CK(clk),
  .Q(\sresult[26][2] ),
  .QN(_05369_)
);

DFF_X1 \sresult[26][3]$_DFFE_PP_  (
  .D(_00315_),
  .CK(clk),
  .Q(\sresult[26][3] ),
  .QN(_05368_)
);

DFF_X1 \sresult[26][4]$_DFFE_PP_  (
  .D(_00316_),
  .CK(clk),
  .Q(\sresult[26][4] ),
  .QN(_05367_)
);

DFF_X1 \sresult[26][5]$_DFFE_PP_  (
  .D(_00317_),
  .CK(clk),
  .Q(\sresult[26][5] ),
  .QN(_05366_)
);

DFF_X1 \sresult[26][6]$_DFFE_PP_  (
  .D(_00318_),
  .CK(clk),
  .Q(\sresult[26][6] ),
  .QN(_05365_)
);

DFF_X1 \sresult[26][7]$_DFFE_PP_  (
  .D(_00319_),
  .CK(clk),
  .Q(\sresult[26][7] ),
  .QN(_05364_)
);

DFF_X1 \sresult[26][8]$_DFFE_PP_  (
  .D(_00320_),
  .CK(clk),
  .Q(\sresult[26][8] ),
  .QN(_05363_)
);

DFF_X1 \sresult[26][9]$_DFFE_PP_  (
  .D(_00321_),
  .CK(clk),
  .Q(\sresult[26][9] ),
  .QN(_05362_)
);

DFF_X1 \sresult[27][0]$_DFFE_PP_  (
  .D(_00324_),
  .CK(clk),
  .Q(\sresult[27][0] ),
  .QN(_05359_)
);

DFF_X1 \sresult[27][10]$_DFFE_PP_  (
  .D(_00334_),
  .CK(clk),
  .Q(\sresult[27][10] ),
  .QN(_05349_)
);

DFF_X1 \sresult[27][11]$_DFFE_PP_  (
  .D(_00335_),
  .CK(clk),
  .Q(\sresult[27][11] ),
  .QN(_05348_)
);

DFF_X1 \sresult[27][1]$_DFFE_PP_  (
  .D(_00325_),
  .CK(clk),
  .Q(\sresult[27][1] ),
  .QN(_05358_)
);

DFF_X1 \sresult[27][2]$_DFFE_PP_  (
  .D(_00326_),
  .CK(clk),
  .Q(\sresult[27][2] ),
  .QN(_05357_)
);

DFF_X1 \sresult[27][3]$_DFFE_PP_  (
  .D(_00327_),
  .CK(clk),
  .Q(\sresult[27][3] ),
  .QN(_05356_)
);

DFF_X1 \sresult[27][4]$_DFFE_PP_  (
  .D(_00328_),
  .CK(clk),
  .Q(\sresult[27][4] ),
  .QN(_05355_)
);

DFF_X1 \sresult[27][5]$_DFFE_PP_  (
  .D(_00329_),
  .CK(clk),
  .Q(\sresult[27][5] ),
  .QN(_05354_)
);

DFF_X1 \sresult[27][6]$_DFFE_PP_  (
  .D(_00330_),
  .CK(clk),
  .Q(\sresult[27][6] ),
  .QN(_05353_)
);

DFF_X1 \sresult[27][7]$_DFFE_PP_  (
  .D(_00331_),
  .CK(clk),
  .Q(\sresult[27][7] ),
  .QN(_05352_)
);

DFF_X1 \sresult[27][8]$_DFFE_PP_  (
  .D(_00332_),
  .CK(clk),
  .Q(\sresult[27][8] ),
  .QN(_05351_)
);

DFF_X1 \sresult[27][9]$_DFFE_PP_  (
  .D(_00333_),
  .CK(clk),
  .Q(\sresult[27][9] ),
  .QN(_05350_)
);

DFF_X1 \sresult[28][0]$_DFFE_PP_  (
  .D(_00336_),
  .CK(clk),
  .Q(\sresult[28][0] ),
  .QN(_05347_)
);

DFF_X1 \sresult[28][10]$_DFFE_PP_  (
  .D(_00346_),
  .CK(clk),
  .Q(\sresult[28][10] ),
  .QN(_05337_)
);

DFF_X1 \sresult[28][11]$_DFFE_PP_  (
  .D(_00347_),
  .CK(clk),
  .Q(\sresult[28][11] ),
  .QN(_05336_)
);

DFF_X1 \sresult[28][1]$_DFFE_PP_  (
  .D(_00337_),
  .CK(clk),
  .Q(\sresult[28][1] ),
  .QN(_05346_)
);

DFF_X1 \sresult[28][2]$_DFFE_PP_  (
  .D(_00338_),
  .CK(clk),
  .Q(\sresult[28][2] ),
  .QN(_05345_)
);

DFF_X1 \sresult[28][3]$_DFFE_PP_  (
  .D(_00339_),
  .CK(clk),
  .Q(\sresult[28][3] ),
  .QN(_05344_)
);

DFF_X1 \sresult[28][4]$_DFFE_PP_  (
  .D(_00340_),
  .CK(clk),
  .Q(\sresult[28][4] ),
  .QN(_05343_)
);

DFF_X1 \sresult[28][5]$_DFFE_PP_  (
  .D(_00341_),
  .CK(clk),
  .Q(\sresult[28][5] ),
  .QN(_05342_)
);

DFF_X1 \sresult[28][6]$_DFFE_PP_  (
  .D(_00342_),
  .CK(clk),
  .Q(\sresult[28][6] ),
  .QN(_05341_)
);

DFF_X1 \sresult[28][7]$_DFFE_PP_  (
  .D(_00343_),
  .CK(clk),
  .Q(\sresult[28][7] ),
  .QN(_05340_)
);

DFF_X1 \sresult[28][8]$_DFFE_PP_  (
  .D(_00344_),
  .CK(clk),
  .Q(\sresult[28][8] ),
  .QN(_05339_)
);

DFF_X1 \sresult[28][9]$_DFFE_PP_  (
  .D(_00345_),
  .CK(clk),
  .Q(\sresult[28][9] ),
  .QN(_05338_)
);

DFF_X1 \sresult[29][0]$_DFFE_PP_  (
  .D(_00348_),
  .CK(clk),
  .Q(\sresult[29][0] ),
  .QN(_05335_)
);

DFF_X1 \sresult[29][10]$_DFFE_PP_  (
  .D(_00358_),
  .CK(clk),
  .Q(\sresult[29][10] ),
  .QN(_05325_)
);

DFF_X1 \sresult[29][11]$_DFFE_PP_  (
  .D(_00359_),
  .CK(clk),
  .Q(\sresult[29][11] ),
  .QN(_05324_)
);

DFF_X1 \sresult[29][1]$_DFFE_PP_  (
  .D(_00349_),
  .CK(clk),
  .Q(\sresult[29][1] ),
  .QN(_05334_)
);

DFF_X1 \sresult[29][2]$_DFFE_PP_  (
  .D(_00350_),
  .CK(clk),
  .Q(\sresult[29][2] ),
  .QN(_05333_)
);

DFF_X1 \sresult[29][3]$_DFFE_PP_  (
  .D(_00351_),
  .CK(clk),
  .Q(\sresult[29][3] ),
  .QN(_05332_)
);

DFF_X1 \sresult[29][4]$_DFFE_PP_  (
  .D(_00352_),
  .CK(clk),
  .Q(\sresult[29][4] ),
  .QN(_05331_)
);

DFF_X1 \sresult[29][5]$_DFFE_PP_  (
  .D(_00353_),
  .CK(clk),
  .Q(\sresult[29][5] ),
  .QN(_05330_)
);

DFF_X1 \sresult[29][6]$_DFFE_PP_  (
  .D(_00354_),
  .CK(clk),
  .Q(\sresult[29][6] ),
  .QN(_05329_)
);

DFF_X1 \sresult[29][7]$_DFFE_PP_  (
  .D(_00355_),
  .CK(clk),
  .Q(\sresult[29][7] ),
  .QN(_05328_)
);

DFF_X1 \sresult[29][8]$_DFFE_PP_  (
  .D(_00356_),
  .CK(clk),
  .Q(\sresult[29][8] ),
  .QN(_05327_)
);

DFF_X1 \sresult[29][9]$_DFFE_PP_  (
  .D(_00357_),
  .CK(clk),
  .Q(\sresult[29][9] ),
  .QN(_05326_)
);

DFF_X1 \sresult[2][0]$_DFFE_PP_  (
  .D(_00024_),
  .CK(clk),
  .Q(\sresult[2][0] ),
  .QN(_05659_)
);

DFF_X1 \sresult[2][10]$_DFFE_PP_  (
  .D(_00034_),
  .CK(clk),
  .Q(\sresult[2][10] ),
  .QN(_05649_)
);

DFF_X1 \sresult[2][11]$_DFFE_PP_  (
  .D(_00035_),
  .CK(clk),
  .Q(\sresult[2][11] ),
  .QN(_05648_)
);

DFF_X1 \sresult[2][1]$_DFFE_PP_  (
  .D(_00025_),
  .CK(clk),
  .Q(\sresult[2][1] ),
  .QN(_05658_)
);

DFF_X1 \sresult[2][2]$_DFFE_PP_  (
  .D(_00026_),
  .CK(clk),
  .Q(\sresult[2][2] ),
  .QN(_05657_)
);

DFF_X1 \sresult[2][3]$_DFFE_PP_  (
  .D(_00027_),
  .CK(clk),
  .Q(\sresult[2][3] ),
  .QN(_05656_)
);

DFF_X1 \sresult[2][4]$_DFFE_PP_  (
  .D(_00028_),
  .CK(clk),
  .Q(\sresult[2][4] ),
  .QN(_05655_)
);

DFF_X1 \sresult[2][5]$_DFFE_PP_  (
  .D(_00029_),
  .CK(clk),
  .Q(\sresult[2][5] ),
  .QN(_05654_)
);

DFF_X1 \sresult[2][6]$_DFFE_PP_  (
  .D(_00030_),
  .CK(clk),
  .Q(\sresult[2][6] ),
  .QN(_05653_)
);

DFF_X1 \sresult[2][7]$_DFFE_PP_  (
  .D(_00031_),
  .CK(clk),
  .Q(\sresult[2][7] ),
  .QN(_05652_)
);

DFF_X1 \sresult[2][8]$_DFFE_PP_  (
  .D(_00032_),
  .CK(clk),
  .Q(\sresult[2][8] ),
  .QN(_05651_)
);

DFF_X1 \sresult[2][9]$_DFFE_PP_  (
  .D(_00033_),
  .CK(clk),
  .Q(\sresult[2][9] ),
  .QN(_05650_)
);

DFF_X1 \sresult[30][0]$_DFFE_PP_  (
  .D(_00360_),
  .CK(clk),
  .Q(\sresult[30][0] ),
  .QN(_05323_)
);

DFF_X1 \sresult[30][10]$_DFFE_PP_  (
  .D(_00370_),
  .CK(clk),
  .Q(\sresult[30][10] ),
  .QN(_05313_)
);

DFF_X1 \sresult[30][11]$_DFFE_PP_  (
  .D(_00371_),
  .CK(clk),
  .Q(\sresult[30][11] ),
  .QN(_05312_)
);

DFF_X1 \sresult[30][1]$_DFFE_PP_  (
  .D(_00361_),
  .CK(clk),
  .Q(\sresult[30][1] ),
  .QN(_05322_)
);

DFF_X1 \sresult[30][2]$_DFFE_PP_  (
  .D(_00362_),
  .CK(clk),
  .Q(\sresult[30][2] ),
  .QN(_05321_)
);

DFF_X1 \sresult[30][3]$_DFFE_PP_  (
  .D(_00363_),
  .CK(clk),
  .Q(\sresult[30][3] ),
  .QN(_05320_)
);

DFF_X1 \sresult[30][4]$_DFFE_PP_  (
  .D(_00364_),
  .CK(clk),
  .Q(\sresult[30][4] ),
  .QN(_05319_)
);

DFF_X1 \sresult[30][5]$_DFFE_PP_  (
  .D(_00365_),
  .CK(clk),
  .Q(\sresult[30][5] ),
  .QN(_05318_)
);

DFF_X1 \sresult[30][6]$_DFFE_PP_  (
  .D(_00366_),
  .CK(clk),
  .Q(\sresult[30][6] ),
  .QN(_05317_)
);

DFF_X1 \sresult[30][7]$_DFFE_PP_  (
  .D(_00367_),
  .CK(clk),
  .Q(\sresult[30][7] ),
  .QN(_05316_)
);

DFF_X1 \sresult[30][8]$_DFFE_PP_  (
  .D(_00368_),
  .CK(clk),
  .Q(\sresult[30][8] ),
  .QN(_05315_)
);

DFF_X1 \sresult[30][9]$_DFFE_PP_  (
  .D(_00369_),
  .CK(clk),
  .Q(\sresult[30][9] ),
  .QN(_05314_)
);

DFF_X1 \sresult[31][0]$_DFFE_PP_  (
  .D(_00372_),
  .CK(clk),
  .Q(\sresult[31][0] ),
  .QN(_05311_)
);

DFF_X1 \sresult[31][10]$_DFFE_PP_  (
  .D(_00382_),
  .CK(clk),
  .Q(\sresult[31][10] ),
  .QN(_05301_)
);

DFF_X1 \sresult[31][11]$_DFFE_PP_  (
  .D(_00383_),
  .CK(clk),
  .Q(\sresult[31][11] ),
  .QN(_05300_)
);

DFF_X1 \sresult[31][1]$_DFFE_PP_  (
  .D(_00373_),
  .CK(clk),
  .Q(\sresult[31][1] ),
  .QN(_05310_)
);

DFF_X1 \sresult[31][2]$_DFFE_PP_  (
  .D(_00374_),
  .CK(clk),
  .Q(\sresult[31][2] ),
  .QN(_05309_)
);

DFF_X1 \sresult[31][3]$_DFFE_PP_  (
  .D(_00375_),
  .CK(clk),
  .Q(\sresult[31][3] ),
  .QN(_05308_)
);

DFF_X1 \sresult[31][4]$_DFFE_PP_  (
  .D(_00376_),
  .CK(clk),
  .Q(\sresult[31][4] ),
  .QN(_05307_)
);

DFF_X1 \sresult[31][5]$_DFFE_PP_  (
  .D(_00377_),
  .CK(clk),
  .Q(\sresult[31][5] ),
  .QN(_05306_)
);

DFF_X1 \sresult[31][6]$_DFFE_PP_  (
  .D(_00378_),
  .CK(clk),
  .Q(\sresult[31][6] ),
  .QN(_05305_)
);

DFF_X1 \sresult[31][7]$_DFFE_PP_  (
  .D(_00379_),
  .CK(clk),
  .Q(\sresult[31][7] ),
  .QN(_05304_)
);

DFF_X1 \sresult[31][8]$_DFFE_PP_  (
  .D(_00380_),
  .CK(clk),
  .Q(\sresult[31][8] ),
  .QN(_05303_)
);

DFF_X1 \sresult[31][9]$_DFFE_PP_  (
  .D(_00381_),
  .CK(clk),
  .Q(\sresult[31][9] ),
  .QN(_05302_)
);

DFF_X1 \sresult[32][0]$_DFFE_PP_  (
  .D(_00384_),
  .CK(clk),
  .Q(\sresult[32][0] ),
  .QN(_05299_)
);

DFF_X1 \sresult[32][10]$_DFFE_PP_  (
  .D(_00394_),
  .CK(clk),
  .Q(\sresult[32][10] ),
  .QN(_05289_)
);

DFF_X1 \sresult[32][11]$_DFFE_PP_  (
  .D(_00395_),
  .CK(clk),
  .Q(\sresult[32][11] ),
  .QN(_05288_)
);

DFF_X1 \sresult[32][1]$_DFFE_PP_  (
  .D(_00385_),
  .CK(clk),
  .Q(\sresult[32][1] ),
  .QN(_05298_)
);

DFF_X1 \sresult[32][2]$_DFFE_PP_  (
  .D(_00386_),
  .CK(clk),
  .Q(\sresult[32][2] ),
  .QN(_05297_)
);

DFF_X1 \sresult[32][3]$_DFFE_PP_  (
  .D(_00387_),
  .CK(clk),
  .Q(\sresult[32][3] ),
  .QN(_05296_)
);

DFF_X1 \sresult[32][4]$_DFFE_PP_  (
  .D(_00388_),
  .CK(clk),
  .Q(\sresult[32][4] ),
  .QN(_05295_)
);

DFF_X1 \sresult[32][5]$_DFFE_PP_  (
  .D(_00389_),
  .CK(clk),
  .Q(\sresult[32][5] ),
  .QN(_05294_)
);

DFF_X1 \sresult[32][6]$_DFFE_PP_  (
  .D(_00390_),
  .CK(clk),
  .Q(\sresult[32][6] ),
  .QN(_05293_)
);

DFF_X1 \sresult[32][7]$_DFFE_PP_  (
  .D(_00391_),
  .CK(clk),
  .Q(\sresult[32][7] ),
  .QN(_05292_)
);

DFF_X1 \sresult[32][8]$_DFFE_PP_  (
  .D(_00392_),
  .CK(clk),
  .Q(\sresult[32][8] ),
  .QN(_05291_)
);

DFF_X1 \sresult[32][9]$_DFFE_PP_  (
  .D(_00393_),
  .CK(clk),
  .Q(\sresult[32][9] ),
  .QN(_05290_)
);

DFF_X1 \sresult[33][0]$_DFFE_PP_  (
  .D(_00396_),
  .CK(clk),
  .Q(\sresult[33][0] ),
  .QN(_05287_)
);

DFF_X1 \sresult[33][10]$_DFFE_PP_  (
  .D(_00406_),
  .CK(clk),
  .Q(\sresult[33][10] ),
  .QN(_05277_)
);

DFF_X1 \sresult[33][11]$_DFFE_PP_  (
  .D(_00407_),
  .CK(clk),
  .Q(\sresult[33][11] ),
  .QN(_05276_)
);

DFF_X1 \sresult[33][1]$_DFFE_PP_  (
  .D(_00397_),
  .CK(clk),
  .Q(\sresult[33][1] ),
  .QN(_05286_)
);

DFF_X1 \sresult[33][2]$_DFFE_PP_  (
  .D(_00398_),
  .CK(clk),
  .Q(\sresult[33][2] ),
  .QN(_05285_)
);

DFF_X1 \sresult[33][3]$_DFFE_PP_  (
  .D(_00399_),
  .CK(clk),
  .Q(\sresult[33][3] ),
  .QN(_05284_)
);

DFF_X1 \sresult[33][4]$_DFFE_PP_  (
  .D(_00400_),
  .CK(clk),
  .Q(\sresult[33][4] ),
  .QN(_05283_)
);

DFF_X1 \sresult[33][5]$_DFFE_PP_  (
  .D(_00401_),
  .CK(clk),
  .Q(\sresult[33][5] ),
  .QN(_05282_)
);

DFF_X1 \sresult[33][6]$_DFFE_PP_  (
  .D(_00402_),
  .CK(clk),
  .Q(\sresult[33][6] ),
  .QN(_05281_)
);

DFF_X1 \sresult[33][7]$_DFFE_PP_  (
  .D(_00403_),
  .CK(clk),
  .Q(\sresult[33][7] ),
  .QN(_05280_)
);

DFF_X1 \sresult[33][8]$_DFFE_PP_  (
  .D(_00404_),
  .CK(clk),
  .Q(\sresult[33][8] ),
  .QN(_05279_)
);

DFF_X1 \sresult[33][9]$_DFFE_PP_  (
  .D(_00405_),
  .CK(clk),
  .Q(\sresult[33][9] ),
  .QN(_05278_)
);

DFF_X1 \sresult[34][0]$_DFFE_PP_  (
  .D(_00408_),
  .CK(clk),
  .Q(\sresult[34][0] ),
  .QN(_05275_)
);

DFF_X1 \sresult[34][10]$_DFFE_PP_  (
  .D(_00418_),
  .CK(clk),
  .Q(\sresult[34][10] ),
  .QN(_05265_)
);

DFF_X1 \sresult[34][11]$_DFFE_PP_  (
  .D(_00419_),
  .CK(clk),
  .Q(\sresult[34][11] ),
  .QN(_05264_)
);

DFF_X1 \sresult[34][1]$_DFFE_PP_  (
  .D(_00409_),
  .CK(clk),
  .Q(\sresult[34][1] ),
  .QN(_05274_)
);

DFF_X1 \sresult[34][2]$_DFFE_PP_  (
  .D(_00410_),
  .CK(clk),
  .Q(\sresult[34][2] ),
  .QN(_05273_)
);

DFF_X1 \sresult[34][3]$_DFFE_PP_  (
  .D(_00411_),
  .CK(clk),
  .Q(\sresult[34][3] ),
  .QN(_05272_)
);

DFF_X1 \sresult[34][4]$_DFFE_PP_  (
  .D(_00412_),
  .CK(clk),
  .Q(\sresult[34][4] ),
  .QN(_05271_)
);

DFF_X1 \sresult[34][5]$_DFFE_PP_  (
  .D(_00413_),
  .CK(clk),
  .Q(\sresult[34][5] ),
  .QN(_05270_)
);

DFF_X1 \sresult[34][6]$_DFFE_PP_  (
  .D(_00414_),
  .CK(clk),
  .Q(\sresult[34][6] ),
  .QN(_05269_)
);

DFF_X1 \sresult[34][7]$_DFFE_PP_  (
  .D(_00415_),
  .CK(clk),
  .Q(\sresult[34][7] ),
  .QN(_05268_)
);

DFF_X1 \sresult[34][8]$_DFFE_PP_  (
  .D(_00416_),
  .CK(clk),
  .Q(\sresult[34][8] ),
  .QN(_05267_)
);

DFF_X1 \sresult[34][9]$_DFFE_PP_  (
  .D(_00417_),
  .CK(clk),
  .Q(\sresult[34][9] ),
  .QN(_05266_)
);

DFF_X1 \sresult[35][0]$_DFFE_PP_  (
  .D(_00420_),
  .CK(clk),
  .Q(\sresult[35][0] ),
  .QN(_05263_)
);

DFF_X1 \sresult[35][10]$_DFFE_PP_  (
  .D(_00430_),
  .CK(clk),
  .Q(\sresult[35][10] ),
  .QN(_05253_)
);

DFF_X1 \sresult[35][11]$_DFFE_PP_  (
  .D(_00431_),
  .CK(clk),
  .Q(\sresult[35][11] ),
  .QN(_05252_)
);

DFF_X1 \sresult[35][1]$_DFFE_PP_  (
  .D(_00421_),
  .CK(clk),
  .Q(\sresult[35][1] ),
  .QN(_05262_)
);

DFF_X1 \sresult[35][2]$_DFFE_PP_  (
  .D(_00422_),
  .CK(clk),
  .Q(\sresult[35][2] ),
  .QN(_05261_)
);

DFF_X1 \sresult[35][3]$_DFFE_PP_  (
  .D(_00423_),
  .CK(clk),
  .Q(\sresult[35][3] ),
  .QN(_05260_)
);

DFF_X1 \sresult[35][4]$_DFFE_PP_  (
  .D(_00424_),
  .CK(clk),
  .Q(\sresult[35][4] ),
  .QN(_05259_)
);

DFF_X1 \sresult[35][5]$_DFFE_PP_  (
  .D(_00425_),
  .CK(clk),
  .Q(\sresult[35][5] ),
  .QN(_05258_)
);

DFF_X1 \sresult[35][6]$_DFFE_PP_  (
  .D(_00426_),
  .CK(clk),
  .Q(\sresult[35][6] ),
  .QN(_05257_)
);

DFF_X1 \sresult[35][7]$_DFFE_PP_  (
  .D(_00427_),
  .CK(clk),
  .Q(\sresult[35][7] ),
  .QN(_05256_)
);

DFF_X1 \sresult[35][8]$_DFFE_PP_  (
  .D(_00428_),
  .CK(clk),
  .Q(\sresult[35][8] ),
  .QN(_05255_)
);

DFF_X1 \sresult[35][9]$_DFFE_PP_  (
  .D(_00429_),
  .CK(clk),
  .Q(\sresult[35][9] ),
  .QN(_05254_)
);

DFF_X1 \sresult[36][0]$_DFFE_PP_  (
  .D(_00432_),
  .CK(clk),
  .Q(\sresult[36][0] ),
  .QN(_05251_)
);

DFF_X1 \sresult[36][10]$_DFFE_PP_  (
  .D(_00442_),
  .CK(clk),
  .Q(\sresult[36][10] ),
  .QN(_05241_)
);

DFF_X1 \sresult[36][11]$_DFFE_PP_  (
  .D(_00443_),
  .CK(clk),
  .Q(\sresult[36][11] ),
  .QN(_05240_)
);

DFF_X1 \sresult[36][1]$_DFFE_PP_  (
  .D(_00433_),
  .CK(clk),
  .Q(\sresult[36][1] ),
  .QN(_05250_)
);

DFF_X1 \sresult[36][2]$_DFFE_PP_  (
  .D(_00434_),
  .CK(clk),
  .Q(\sresult[36][2] ),
  .QN(_05249_)
);

DFF_X1 \sresult[36][3]$_DFFE_PP_  (
  .D(_00435_),
  .CK(clk),
  .Q(\sresult[36][3] ),
  .QN(_05248_)
);

DFF_X1 \sresult[36][4]$_DFFE_PP_  (
  .D(_00436_),
  .CK(clk),
  .Q(\sresult[36][4] ),
  .QN(_05247_)
);

DFF_X1 \sresult[36][5]$_DFFE_PP_  (
  .D(_00437_),
  .CK(clk),
  .Q(\sresult[36][5] ),
  .QN(_05246_)
);

DFF_X1 \sresult[36][6]$_DFFE_PP_  (
  .D(_00438_),
  .CK(clk),
  .Q(\sresult[36][6] ),
  .QN(_05245_)
);

DFF_X1 \sresult[36][7]$_DFFE_PP_  (
  .D(_00439_),
  .CK(clk),
  .Q(\sresult[36][7] ),
  .QN(_05244_)
);

DFF_X1 \sresult[36][8]$_DFFE_PP_  (
  .D(_00440_),
  .CK(clk),
  .Q(\sresult[36][8] ),
  .QN(_05243_)
);

DFF_X1 \sresult[36][9]$_DFFE_PP_  (
  .D(_00441_),
  .CK(clk),
  .Q(\sresult[36][9] ),
  .QN(_05242_)
);

DFF_X1 \sresult[37][0]$_DFFE_PP_  (
  .D(_00444_),
  .CK(clk),
  .Q(\sresult[37][0] ),
  .QN(_05239_)
);

DFF_X1 \sresult[37][10]$_DFFE_PP_  (
  .D(_00454_),
  .CK(clk),
  .Q(\sresult[37][10] ),
  .QN(_05229_)
);

DFF_X1 \sresult[37][11]$_DFFE_PP_  (
  .D(_00455_),
  .CK(clk),
  .Q(\sresult[37][11] ),
  .QN(_05228_)
);

DFF_X1 \sresult[37][1]$_DFFE_PP_  (
  .D(_00445_),
  .CK(clk),
  .Q(\sresult[37][1] ),
  .QN(_05238_)
);

DFF_X1 \sresult[37][2]$_DFFE_PP_  (
  .D(_00446_),
  .CK(clk),
  .Q(\sresult[37][2] ),
  .QN(_05237_)
);

DFF_X1 \sresult[37][3]$_DFFE_PP_  (
  .D(_00447_),
  .CK(clk),
  .Q(\sresult[37][3] ),
  .QN(_05236_)
);

DFF_X1 \sresult[37][4]$_DFFE_PP_  (
  .D(_00448_),
  .CK(clk),
  .Q(\sresult[37][4] ),
  .QN(_05235_)
);

DFF_X1 \sresult[37][5]$_DFFE_PP_  (
  .D(_00449_),
  .CK(clk),
  .Q(\sresult[37][5] ),
  .QN(_05234_)
);

DFF_X1 \sresult[37][6]$_DFFE_PP_  (
  .D(_00450_),
  .CK(clk),
  .Q(\sresult[37][6] ),
  .QN(_05233_)
);

DFF_X1 \sresult[37][7]$_DFFE_PP_  (
  .D(_00451_),
  .CK(clk),
  .Q(\sresult[37][7] ),
  .QN(_05232_)
);

DFF_X1 \sresult[37][8]$_DFFE_PP_  (
  .D(_00452_),
  .CK(clk),
  .Q(\sresult[37][8] ),
  .QN(_05231_)
);

DFF_X1 \sresult[37][9]$_DFFE_PP_  (
  .D(_00453_),
  .CK(clk),
  .Q(\sresult[37][9] ),
  .QN(_05230_)
);

DFF_X1 \sresult[38][0]$_DFFE_PP_  (
  .D(_00456_),
  .CK(clk),
  .Q(\sresult[38][0] ),
  .QN(_05227_)
);

DFF_X1 \sresult[38][10]$_DFFE_PP_  (
  .D(_00466_),
  .CK(clk),
  .Q(\sresult[38][10] ),
  .QN(_05217_)
);

DFF_X1 \sresult[38][11]$_DFFE_PP_  (
  .D(_00467_),
  .CK(clk),
  .Q(\sresult[38][11] ),
  .QN(_05216_)
);

DFF_X1 \sresult[38][1]$_DFFE_PP_  (
  .D(_00457_),
  .CK(clk),
  .Q(\sresult[38][1] ),
  .QN(_05226_)
);

DFF_X1 \sresult[38][2]$_DFFE_PP_  (
  .D(_00458_),
  .CK(clk),
  .Q(\sresult[38][2] ),
  .QN(_05225_)
);

DFF_X1 \sresult[38][3]$_DFFE_PP_  (
  .D(_00459_),
  .CK(clk),
  .Q(\sresult[38][3] ),
  .QN(_05224_)
);

DFF_X1 \sresult[38][4]$_DFFE_PP_  (
  .D(_00460_),
  .CK(clk),
  .Q(\sresult[38][4] ),
  .QN(_05223_)
);

DFF_X1 \sresult[38][5]$_DFFE_PP_  (
  .D(_00461_),
  .CK(clk),
  .Q(\sresult[38][5] ),
  .QN(_05222_)
);

DFF_X1 \sresult[38][6]$_DFFE_PP_  (
  .D(_00462_),
  .CK(clk),
  .Q(\sresult[38][6] ),
  .QN(_05221_)
);

DFF_X1 \sresult[38][7]$_DFFE_PP_  (
  .D(_00463_),
  .CK(clk),
  .Q(\sresult[38][7] ),
  .QN(_05220_)
);

DFF_X1 \sresult[38][8]$_DFFE_PP_  (
  .D(_00464_),
  .CK(clk),
  .Q(\sresult[38][8] ),
  .QN(_05219_)
);

DFF_X1 \sresult[38][9]$_DFFE_PP_  (
  .D(_00465_),
  .CK(clk),
  .Q(\sresult[38][9] ),
  .QN(_05218_)
);

DFF_X1 \sresult[39][0]$_DFFE_PP_  (
  .D(_00468_),
  .CK(clk),
  .Q(\sresult[39][0] ),
  .QN(_05215_)
);

DFF_X1 \sresult[39][10]$_DFFE_PP_  (
  .D(_00478_),
  .CK(clk),
  .Q(\sresult[39][10] ),
  .QN(_05205_)
);

DFF_X1 \sresult[39][11]$_DFFE_PP_  (
  .D(_00479_),
  .CK(clk),
  .Q(\sresult[39][11] ),
  .QN(_05204_)
);

DFF_X1 \sresult[39][1]$_DFFE_PP_  (
  .D(_00469_),
  .CK(clk),
  .Q(\sresult[39][1] ),
  .QN(_05214_)
);

DFF_X1 \sresult[39][2]$_DFFE_PP_  (
  .D(_00470_),
  .CK(clk),
  .Q(\sresult[39][2] ),
  .QN(_05213_)
);

DFF_X1 \sresult[39][3]$_DFFE_PP_  (
  .D(_00471_),
  .CK(clk),
  .Q(\sresult[39][3] ),
  .QN(_05212_)
);

DFF_X1 \sresult[39][4]$_DFFE_PP_  (
  .D(_00472_),
  .CK(clk),
  .Q(\sresult[39][4] ),
  .QN(_05211_)
);

DFF_X1 \sresult[39][5]$_DFFE_PP_  (
  .D(_00473_),
  .CK(clk),
  .Q(\sresult[39][5] ),
  .QN(_05210_)
);

DFF_X1 \sresult[39][6]$_DFFE_PP_  (
  .D(_00474_),
  .CK(clk),
  .Q(\sresult[39][6] ),
  .QN(_05209_)
);

DFF_X1 \sresult[39][7]$_DFFE_PP_  (
  .D(_00475_),
  .CK(clk),
  .Q(\sresult[39][7] ),
  .QN(_05208_)
);

DFF_X1 \sresult[39][8]$_DFFE_PP_  (
  .D(_00476_),
  .CK(clk),
  .Q(\sresult[39][8] ),
  .QN(_05207_)
);

DFF_X1 \sresult[39][9]$_DFFE_PP_  (
  .D(_00477_),
  .CK(clk),
  .Q(\sresult[39][9] ),
  .QN(_05206_)
);

DFF_X1 \sresult[3][0]$_DFFE_PP_  (
  .D(_00036_),
  .CK(clk),
  .Q(\sresult[3][0] ),
  .QN(_05647_)
);

DFF_X1 \sresult[3][10]$_DFFE_PP_  (
  .D(_00046_),
  .CK(clk),
  .Q(\sresult[3][10] ),
  .QN(_05637_)
);

DFF_X1 \sresult[3][11]$_DFFE_PP_  (
  .D(_00047_),
  .CK(clk),
  .Q(\sresult[3][11] ),
  .QN(_05636_)
);

DFF_X1 \sresult[3][1]$_DFFE_PP_  (
  .D(_00037_),
  .CK(clk),
  .Q(\sresult[3][1] ),
  .QN(_05646_)
);

DFF_X1 \sresult[3][2]$_DFFE_PP_  (
  .D(_00038_),
  .CK(clk),
  .Q(\sresult[3][2] ),
  .QN(_05645_)
);

DFF_X1 \sresult[3][3]$_DFFE_PP_  (
  .D(_00039_),
  .CK(clk),
  .Q(\sresult[3][3] ),
  .QN(_05644_)
);

DFF_X1 \sresult[3][4]$_DFFE_PP_  (
  .D(_00040_),
  .CK(clk),
  .Q(\sresult[3][4] ),
  .QN(_05643_)
);

DFF_X1 \sresult[3][5]$_DFFE_PP_  (
  .D(_00041_),
  .CK(clk),
  .Q(\sresult[3][5] ),
  .QN(_05642_)
);

DFF_X1 \sresult[3][6]$_DFFE_PP_  (
  .D(_00042_),
  .CK(clk),
  .Q(\sresult[3][6] ),
  .QN(_05641_)
);

DFF_X1 \sresult[3][7]$_DFFE_PP_  (
  .D(_00043_),
  .CK(clk),
  .Q(\sresult[3][7] ),
  .QN(_05640_)
);

DFF_X1 \sresult[3][8]$_DFFE_PP_  (
  .D(_00044_),
  .CK(clk),
  .Q(\sresult[3][8] ),
  .QN(_05639_)
);

DFF_X1 \sresult[3][9]$_DFFE_PP_  (
  .D(_00045_),
  .CK(clk),
  .Q(\sresult[3][9] ),
  .QN(_05638_)
);

DFF_X1 \sresult[40][0]$_DFFE_PP_  (
  .D(_00480_),
  .CK(clk),
  .Q(\sresult[40][0] ),
  .QN(_05203_)
);

DFF_X1 \sresult[40][10]$_DFFE_PP_  (
  .D(_00490_),
  .CK(clk),
  .Q(\sresult[40][10] ),
  .QN(_05193_)
);

DFF_X1 \sresult[40][11]$_DFFE_PP_  (
  .D(_00491_),
  .CK(clk),
  .Q(\sresult[40][11] ),
  .QN(_05192_)
);

DFF_X1 \sresult[40][1]$_DFFE_PP_  (
  .D(_00481_),
  .CK(clk),
  .Q(\sresult[40][1] ),
  .QN(_05202_)
);

DFF_X1 \sresult[40][2]$_DFFE_PP_  (
  .D(_00482_),
  .CK(clk),
  .Q(\sresult[40][2] ),
  .QN(_05201_)
);

DFF_X1 \sresult[40][3]$_DFFE_PP_  (
  .D(_00483_),
  .CK(clk),
  .Q(\sresult[40][3] ),
  .QN(_05200_)
);

DFF_X1 \sresult[40][4]$_DFFE_PP_  (
  .D(_00484_),
  .CK(clk),
  .Q(\sresult[40][4] ),
  .QN(_05199_)
);

DFF_X1 \sresult[40][5]$_DFFE_PP_  (
  .D(_00485_),
  .CK(clk),
  .Q(\sresult[40][5] ),
  .QN(_05198_)
);

DFF_X1 \sresult[40][6]$_DFFE_PP_  (
  .D(_00486_),
  .CK(clk),
  .Q(\sresult[40][6] ),
  .QN(_05197_)
);

DFF_X1 \sresult[40][7]$_DFFE_PP_  (
  .D(_00487_),
  .CK(clk),
  .Q(\sresult[40][7] ),
  .QN(_05196_)
);

DFF_X1 \sresult[40][8]$_DFFE_PP_  (
  .D(_00488_),
  .CK(clk),
  .Q(\sresult[40][8] ),
  .QN(_05195_)
);

DFF_X1 \sresult[40][9]$_DFFE_PP_  (
  .D(_00489_),
  .CK(clk),
  .Q(\sresult[40][9] ),
  .QN(_05194_)
);

DFF_X1 \sresult[41][0]$_DFFE_PP_  (
  .D(_00492_),
  .CK(clk),
  .Q(\sresult[41][0] ),
  .QN(_05191_)
);

DFF_X1 \sresult[41][10]$_DFFE_PP_  (
  .D(_00502_),
  .CK(clk),
  .Q(\sresult[41][10] ),
  .QN(_05181_)
);

DFF_X1 \sresult[41][11]$_DFFE_PP_  (
  .D(_00503_),
  .CK(clk),
  .Q(\sresult[41][11] ),
  .QN(_05180_)
);

DFF_X1 \sresult[41][1]$_DFFE_PP_  (
  .D(_00493_),
  .CK(clk),
  .Q(\sresult[41][1] ),
  .QN(_05190_)
);

DFF_X1 \sresult[41][2]$_DFFE_PP_  (
  .D(_00494_),
  .CK(clk),
  .Q(\sresult[41][2] ),
  .QN(_05189_)
);

DFF_X1 \sresult[41][3]$_DFFE_PP_  (
  .D(_00495_),
  .CK(clk),
  .Q(\sresult[41][3] ),
  .QN(_05188_)
);

DFF_X1 \sresult[41][4]$_DFFE_PP_  (
  .D(_00496_),
  .CK(clk),
  .Q(\sresult[41][4] ),
  .QN(_05187_)
);

DFF_X1 \sresult[41][5]$_DFFE_PP_  (
  .D(_00497_),
  .CK(clk),
  .Q(\sresult[41][5] ),
  .QN(_05186_)
);

DFF_X1 \sresult[41][6]$_DFFE_PP_  (
  .D(_00498_),
  .CK(clk),
  .Q(\sresult[41][6] ),
  .QN(_05185_)
);

DFF_X1 \sresult[41][7]$_DFFE_PP_  (
  .D(_00499_),
  .CK(clk),
  .Q(\sresult[41][7] ),
  .QN(_05184_)
);

DFF_X1 \sresult[41][8]$_DFFE_PP_  (
  .D(_00500_),
  .CK(clk),
  .Q(\sresult[41][8] ),
  .QN(_05183_)
);

DFF_X1 \sresult[41][9]$_DFFE_PP_  (
  .D(_00501_),
  .CK(clk),
  .Q(\sresult[41][9] ),
  .QN(_05182_)
);

DFF_X1 \sresult[42][0]$_DFFE_PP_  (
  .D(_00504_),
  .CK(clk),
  .Q(\sresult[42][0] ),
  .QN(_05179_)
);

DFF_X1 \sresult[42][10]$_DFFE_PP_  (
  .D(_00514_),
  .CK(clk),
  .Q(\sresult[42][10] ),
  .QN(_05169_)
);

DFF_X1 \sresult[42][11]$_DFFE_PP_  (
  .D(_00515_),
  .CK(clk),
  .Q(\sresult[42][11] ),
  .QN(_05168_)
);

DFF_X1 \sresult[42][1]$_DFFE_PP_  (
  .D(_00505_),
  .CK(clk),
  .Q(\sresult[42][1] ),
  .QN(_05178_)
);

DFF_X1 \sresult[42][2]$_DFFE_PP_  (
  .D(_00506_),
  .CK(clk),
  .Q(\sresult[42][2] ),
  .QN(_05177_)
);

DFF_X1 \sresult[42][3]$_DFFE_PP_  (
  .D(_00507_),
  .CK(clk),
  .Q(\sresult[42][3] ),
  .QN(_05176_)
);

DFF_X1 \sresult[42][4]$_DFFE_PP_  (
  .D(_00508_),
  .CK(clk),
  .Q(\sresult[42][4] ),
  .QN(_05175_)
);

DFF_X1 \sresult[42][5]$_DFFE_PP_  (
  .D(_00509_),
  .CK(clk),
  .Q(\sresult[42][5] ),
  .QN(_05174_)
);

DFF_X1 \sresult[42][6]$_DFFE_PP_  (
  .D(_00510_),
  .CK(clk),
  .Q(\sresult[42][6] ),
  .QN(_05173_)
);

DFF_X1 \sresult[42][7]$_DFFE_PP_  (
  .D(_00511_),
  .CK(clk),
  .Q(\sresult[42][7] ),
  .QN(_05172_)
);

DFF_X1 \sresult[42][8]$_DFFE_PP_  (
  .D(_00512_),
  .CK(clk),
  .Q(\sresult[42][8] ),
  .QN(_05171_)
);

DFF_X1 \sresult[42][9]$_DFFE_PP_  (
  .D(_00513_),
  .CK(clk),
  .Q(\sresult[42][9] ),
  .QN(_05170_)
);

DFF_X1 \sresult[43][0]$_DFFE_PP_  (
  .D(_00516_),
  .CK(clk),
  .Q(\sresult[43][0] ),
  .QN(_05167_)
);

DFF_X1 \sresult[43][10]$_DFFE_PP_  (
  .D(_00526_),
  .CK(clk),
  .Q(\sresult[43][10] ),
  .QN(_05157_)
);

DFF_X1 \sresult[43][11]$_DFFE_PP_  (
  .D(_00527_),
  .CK(clk),
  .Q(\sresult[43][11] ),
  .QN(_05156_)
);

DFF_X1 \sresult[43][1]$_DFFE_PP_  (
  .D(_00517_),
  .CK(clk),
  .Q(\sresult[43][1] ),
  .QN(_05166_)
);

DFF_X1 \sresult[43][2]$_DFFE_PP_  (
  .D(_00518_),
  .CK(clk),
  .Q(\sresult[43][2] ),
  .QN(_05165_)
);

DFF_X1 \sresult[43][3]$_DFFE_PP_  (
  .D(_00519_),
  .CK(clk),
  .Q(\sresult[43][3] ),
  .QN(_05164_)
);

DFF_X1 \sresult[43][4]$_DFFE_PP_  (
  .D(_00520_),
  .CK(clk),
  .Q(\sresult[43][4] ),
  .QN(_05163_)
);

DFF_X1 \sresult[43][5]$_DFFE_PP_  (
  .D(_00521_),
  .CK(clk),
  .Q(\sresult[43][5] ),
  .QN(_05162_)
);

DFF_X1 \sresult[43][6]$_DFFE_PP_  (
  .D(_00522_),
  .CK(clk),
  .Q(\sresult[43][6] ),
  .QN(_05161_)
);

DFF_X1 \sresult[43][7]$_DFFE_PP_  (
  .D(_00523_),
  .CK(clk),
  .Q(\sresult[43][7] ),
  .QN(_05160_)
);

DFF_X1 \sresult[43][8]$_DFFE_PP_  (
  .D(_00524_),
  .CK(clk),
  .Q(\sresult[43][8] ),
  .QN(_05159_)
);

DFF_X1 \sresult[43][9]$_DFFE_PP_  (
  .D(_00525_),
  .CK(clk),
  .Q(\sresult[43][9] ),
  .QN(_05158_)
);

DFF_X1 \sresult[44][0]$_DFFE_PP_  (
  .D(_00528_),
  .CK(clk),
  .Q(\sresult[44][0] ),
  .QN(_05155_)
);

DFF_X1 \sresult[44][10]$_DFFE_PP_  (
  .D(_00538_),
  .CK(clk),
  .Q(\sresult[44][10] ),
  .QN(_05145_)
);

DFF_X1 \sresult[44][11]$_DFFE_PP_  (
  .D(_00539_),
  .CK(clk),
  .Q(\sresult[44][11] ),
  .QN(_05144_)
);

DFF_X1 \sresult[44][1]$_DFFE_PP_  (
  .D(_00529_),
  .CK(clk),
  .Q(\sresult[44][1] ),
  .QN(_05154_)
);

DFF_X1 \sresult[44][2]$_DFFE_PP_  (
  .D(_00530_),
  .CK(clk),
  .Q(\sresult[44][2] ),
  .QN(_05153_)
);

DFF_X1 \sresult[44][3]$_DFFE_PP_  (
  .D(_00531_),
  .CK(clk),
  .Q(\sresult[44][3] ),
  .QN(_05152_)
);

DFF_X1 \sresult[44][4]$_DFFE_PP_  (
  .D(_00532_),
  .CK(clk),
  .Q(\sresult[44][4] ),
  .QN(_05151_)
);

DFF_X1 \sresult[44][5]$_DFFE_PP_  (
  .D(_00533_),
  .CK(clk),
  .Q(\sresult[44][5] ),
  .QN(_05150_)
);

DFF_X1 \sresult[44][6]$_DFFE_PP_  (
  .D(_00534_),
  .CK(clk),
  .Q(\sresult[44][6] ),
  .QN(_05149_)
);

DFF_X1 \sresult[44][7]$_DFFE_PP_  (
  .D(_00535_),
  .CK(clk),
  .Q(\sresult[44][7] ),
  .QN(_05148_)
);

DFF_X1 \sresult[44][8]$_DFFE_PP_  (
  .D(_00536_),
  .CK(clk),
  .Q(\sresult[44][8] ),
  .QN(_05147_)
);

DFF_X1 \sresult[44][9]$_DFFE_PP_  (
  .D(_00537_),
  .CK(clk),
  .Q(\sresult[44][9] ),
  .QN(_05146_)
);

DFF_X1 \sresult[45][0]$_DFFE_PP_  (
  .D(_00540_),
  .CK(clk),
  .Q(\sresult[45][0] ),
  .QN(_05143_)
);

DFF_X1 \sresult[45][10]$_DFFE_PP_  (
  .D(_00550_),
  .CK(clk),
  .Q(\sresult[45][10] ),
  .QN(_05133_)
);

DFF_X1 \sresult[45][11]$_DFFE_PP_  (
  .D(_00551_),
  .CK(clk),
  .Q(\sresult[45][11] ),
  .QN(_05132_)
);

DFF_X1 \sresult[45][1]$_DFFE_PP_  (
  .D(_00541_),
  .CK(clk),
  .Q(\sresult[45][1] ),
  .QN(_05142_)
);

DFF_X1 \sresult[45][2]$_DFFE_PP_  (
  .D(_00542_),
  .CK(clk),
  .Q(\sresult[45][2] ),
  .QN(_05141_)
);

DFF_X1 \sresult[45][3]$_DFFE_PP_  (
  .D(_00543_),
  .CK(clk),
  .Q(\sresult[45][3] ),
  .QN(_05140_)
);

DFF_X1 \sresult[45][4]$_DFFE_PP_  (
  .D(_00544_),
  .CK(clk),
  .Q(\sresult[45][4] ),
  .QN(_05139_)
);

DFF_X1 \sresult[45][5]$_DFFE_PP_  (
  .D(_00545_),
  .CK(clk),
  .Q(\sresult[45][5] ),
  .QN(_05138_)
);

DFF_X1 \sresult[45][6]$_DFFE_PP_  (
  .D(_00546_),
  .CK(clk),
  .Q(\sresult[45][6] ),
  .QN(_05137_)
);

DFF_X1 \sresult[45][7]$_DFFE_PP_  (
  .D(_00547_),
  .CK(clk),
  .Q(\sresult[45][7] ),
  .QN(_05136_)
);

DFF_X1 \sresult[45][8]$_DFFE_PP_  (
  .D(_00548_),
  .CK(clk),
  .Q(\sresult[45][8] ),
  .QN(_05135_)
);

DFF_X1 \sresult[45][9]$_DFFE_PP_  (
  .D(_00549_),
  .CK(clk),
  .Q(\sresult[45][9] ),
  .QN(_05134_)
);

DFF_X1 \sresult[46][0]$_DFFE_PP_  (
  .D(_00552_),
  .CK(clk),
  .Q(\sresult[46][0] ),
  .QN(_05131_)
);

DFF_X1 \sresult[46][10]$_DFFE_PP_  (
  .D(_00562_),
  .CK(clk),
  .Q(\sresult[46][10] ),
  .QN(_05121_)
);

DFF_X1 \sresult[46][11]$_DFFE_PP_  (
  .D(_00563_),
  .CK(clk),
  .Q(\sresult[46][11] ),
  .QN(_05120_)
);

DFF_X1 \sresult[46][1]$_DFFE_PP_  (
  .D(_00553_),
  .CK(clk),
  .Q(\sresult[46][1] ),
  .QN(_05130_)
);

DFF_X1 \sresult[46][2]$_DFFE_PP_  (
  .D(_00554_),
  .CK(clk),
  .Q(\sresult[46][2] ),
  .QN(_05129_)
);

DFF_X1 \sresult[46][3]$_DFFE_PP_  (
  .D(_00555_),
  .CK(clk),
  .Q(\sresult[46][3] ),
  .QN(_05128_)
);

DFF_X1 \sresult[46][4]$_DFFE_PP_  (
  .D(_00556_),
  .CK(clk),
  .Q(\sresult[46][4] ),
  .QN(_05127_)
);

DFF_X1 \sresult[46][5]$_DFFE_PP_  (
  .D(_00557_),
  .CK(clk),
  .Q(\sresult[46][5] ),
  .QN(_05126_)
);

DFF_X1 \sresult[46][6]$_DFFE_PP_  (
  .D(_00558_),
  .CK(clk),
  .Q(\sresult[46][6] ),
  .QN(_05125_)
);

DFF_X1 \sresult[46][7]$_DFFE_PP_  (
  .D(_00559_),
  .CK(clk),
  .Q(\sresult[46][7] ),
  .QN(_05124_)
);

DFF_X1 \sresult[46][8]$_DFFE_PP_  (
  .D(_00560_),
  .CK(clk),
  .Q(\sresult[46][8] ),
  .QN(_05123_)
);

DFF_X1 \sresult[46][9]$_DFFE_PP_  (
  .D(_00561_),
  .CK(clk),
  .Q(\sresult[46][9] ),
  .QN(_05122_)
);

DFF_X1 \sresult[47][0]$_DFFE_PP_  (
  .D(_00564_),
  .CK(clk),
  .Q(\sresult[47][0] ),
  .QN(_05119_)
);

DFF_X1 \sresult[47][10]$_DFFE_PP_  (
  .D(_00574_),
  .CK(clk),
  .Q(\sresult[47][10] ),
  .QN(_05109_)
);

DFF_X1 \sresult[47][11]$_DFFE_PP_  (
  .D(_00575_),
  .CK(clk),
  .Q(\sresult[47][11] ),
  .QN(_05108_)
);

DFF_X1 \sresult[47][1]$_DFFE_PP_  (
  .D(_00565_),
  .CK(clk),
  .Q(\sresult[47][1] ),
  .QN(_05118_)
);

DFF_X1 \sresult[47][2]$_DFFE_PP_  (
  .D(_00566_),
  .CK(clk),
  .Q(\sresult[47][2] ),
  .QN(_05117_)
);

DFF_X1 \sresult[47][3]$_DFFE_PP_  (
  .D(_00567_),
  .CK(clk),
  .Q(\sresult[47][3] ),
  .QN(_05116_)
);

DFF_X1 \sresult[47][4]$_DFFE_PP_  (
  .D(_00568_),
  .CK(clk),
  .Q(\sresult[47][4] ),
  .QN(_05115_)
);

DFF_X1 \sresult[47][5]$_DFFE_PP_  (
  .D(_00569_),
  .CK(clk),
  .Q(\sresult[47][5] ),
  .QN(_05114_)
);

DFF_X1 \sresult[47][6]$_DFFE_PP_  (
  .D(_00570_),
  .CK(clk),
  .Q(\sresult[47][6] ),
  .QN(_05113_)
);

DFF_X1 \sresult[47][7]$_DFFE_PP_  (
  .D(_00571_),
  .CK(clk),
  .Q(\sresult[47][7] ),
  .QN(_05112_)
);

DFF_X1 \sresult[47][8]$_DFFE_PP_  (
  .D(_00572_),
  .CK(clk),
  .Q(\sresult[47][8] ),
  .QN(_05111_)
);

DFF_X1 \sresult[47][9]$_DFFE_PP_  (
  .D(_00573_),
  .CK(clk),
  .Q(\sresult[47][9] ),
  .QN(_05110_)
);

DFF_X1 \sresult[48][0]$_DFFE_PP_  (
  .D(_00576_),
  .CK(clk),
  .Q(\sresult[48][0] ),
  .QN(_05107_)
);

DFF_X1 \sresult[48][10]$_DFFE_PP_  (
  .D(_00586_),
  .CK(clk),
  .Q(\sresult[48][10] ),
  .QN(_05097_)
);

DFF_X1 \sresult[48][11]$_DFFE_PP_  (
  .D(_00587_),
  .CK(clk),
  .Q(\sresult[48][11] ),
  .QN(_05096_)
);

DFF_X1 \sresult[48][1]$_DFFE_PP_  (
  .D(_00577_),
  .CK(clk),
  .Q(\sresult[48][1] ),
  .QN(_05106_)
);

DFF_X1 \sresult[48][2]$_DFFE_PP_  (
  .D(_00578_),
  .CK(clk),
  .Q(\sresult[48][2] ),
  .QN(_05105_)
);

DFF_X1 \sresult[48][3]$_DFFE_PP_  (
  .D(_00579_),
  .CK(clk),
  .Q(\sresult[48][3] ),
  .QN(_05104_)
);

DFF_X1 \sresult[48][4]$_DFFE_PP_  (
  .D(_00580_),
  .CK(clk),
  .Q(\sresult[48][4] ),
  .QN(_05103_)
);

DFF_X1 \sresult[48][5]$_DFFE_PP_  (
  .D(_00581_),
  .CK(clk),
  .Q(\sresult[48][5] ),
  .QN(_05102_)
);

DFF_X1 \sresult[48][6]$_DFFE_PP_  (
  .D(_00582_),
  .CK(clk),
  .Q(\sresult[48][6] ),
  .QN(_05101_)
);

DFF_X1 \sresult[48][7]$_DFFE_PP_  (
  .D(_00583_),
  .CK(clk),
  .Q(\sresult[48][7] ),
  .QN(_05100_)
);

DFF_X1 \sresult[48][8]$_DFFE_PP_  (
  .D(_00584_),
  .CK(clk),
  .Q(\sresult[48][8] ),
  .QN(_05099_)
);

DFF_X1 \sresult[48][9]$_DFFE_PP_  (
  .D(_00585_),
  .CK(clk),
  .Q(\sresult[48][9] ),
  .QN(_05098_)
);

DFF_X1 \sresult[49][0]$_DFFE_PP_  (
  .D(_00588_),
  .CK(clk),
  .Q(\sresult[49][0] ),
  .QN(_05095_)
);

DFF_X1 \sresult[49][10]$_DFFE_PP_  (
  .D(_00598_),
  .CK(clk),
  .Q(\sresult[49][10] ),
  .QN(_05085_)
);

DFF_X1 \sresult[49][11]$_DFFE_PP_  (
  .D(_00599_),
  .CK(clk),
  .Q(\sresult[49][11] ),
  .QN(_05084_)
);

DFF_X1 \sresult[49][1]$_DFFE_PP_  (
  .D(_00589_),
  .CK(clk),
  .Q(\sresult[49][1] ),
  .QN(_05094_)
);

DFF_X1 \sresult[49][2]$_DFFE_PP_  (
  .D(_00590_),
  .CK(clk),
  .Q(\sresult[49][2] ),
  .QN(_05093_)
);

DFF_X1 \sresult[49][3]$_DFFE_PP_  (
  .D(_00591_),
  .CK(clk),
  .Q(\sresult[49][3] ),
  .QN(_05092_)
);

DFF_X1 \sresult[49][4]$_DFFE_PP_  (
  .D(_00592_),
  .CK(clk),
  .Q(\sresult[49][4] ),
  .QN(_05091_)
);

DFF_X1 \sresult[49][5]$_DFFE_PP_  (
  .D(_00593_),
  .CK(clk),
  .Q(\sresult[49][5] ),
  .QN(_05090_)
);

DFF_X1 \sresult[49][6]$_DFFE_PP_  (
  .D(_00594_),
  .CK(clk),
  .Q(\sresult[49][6] ),
  .QN(_05089_)
);

DFF_X1 \sresult[49][7]$_DFFE_PP_  (
  .D(_00595_),
  .CK(clk),
  .Q(\sresult[49][7] ),
  .QN(_05088_)
);

DFF_X1 \sresult[49][8]$_DFFE_PP_  (
  .D(_00596_),
  .CK(clk),
  .Q(\sresult[49][8] ),
  .QN(_05087_)
);

DFF_X1 \sresult[49][9]$_DFFE_PP_  (
  .D(_00597_),
  .CK(clk),
  .Q(\sresult[49][9] ),
  .QN(_05086_)
);

DFF_X1 \sresult[4][0]$_DFFE_PP_  (
  .D(_00048_),
  .CK(clk),
  .Q(\sresult[4][0] ),
  .QN(_05635_)
);

DFF_X1 \sresult[4][10]$_DFFE_PP_  (
  .D(_00058_),
  .CK(clk),
  .Q(\sresult[4][10] ),
  .QN(_05625_)
);

DFF_X1 \sresult[4][11]$_DFFE_PP_  (
  .D(_00059_),
  .CK(clk),
  .Q(\sresult[4][11] ),
  .QN(_05624_)
);

DFF_X1 \sresult[4][1]$_DFFE_PP_  (
  .D(_00049_),
  .CK(clk),
  .Q(\sresult[4][1] ),
  .QN(_05634_)
);

DFF_X1 \sresult[4][2]$_DFFE_PP_  (
  .D(_00050_),
  .CK(clk),
  .Q(\sresult[4][2] ),
  .QN(_05633_)
);

DFF_X1 \sresult[4][3]$_DFFE_PP_  (
  .D(_00051_),
  .CK(clk),
  .Q(\sresult[4][3] ),
  .QN(_05632_)
);

DFF_X1 \sresult[4][4]$_DFFE_PP_  (
  .D(_00052_),
  .CK(clk),
  .Q(\sresult[4][4] ),
  .QN(_05631_)
);

DFF_X1 \sresult[4][5]$_DFFE_PP_  (
  .D(_00053_),
  .CK(clk),
  .Q(\sresult[4][5] ),
  .QN(_05630_)
);

DFF_X1 \sresult[4][6]$_DFFE_PP_  (
  .D(_00054_),
  .CK(clk),
  .Q(\sresult[4][6] ),
  .QN(_05629_)
);

DFF_X1 \sresult[4][7]$_DFFE_PP_  (
  .D(_00055_),
  .CK(clk),
  .Q(\sresult[4][7] ),
  .QN(_05628_)
);

DFF_X1 \sresult[4][8]$_DFFE_PP_  (
  .D(_00056_),
  .CK(clk),
  .Q(\sresult[4][8] ),
  .QN(_05627_)
);

DFF_X1 \sresult[4][9]$_DFFE_PP_  (
  .D(_00057_),
  .CK(clk),
  .Q(\sresult[4][9] ),
  .QN(_05626_)
);

DFF_X1 \sresult[50][0]$_DFFE_PP_  (
  .D(_00600_),
  .CK(clk),
  .Q(\sresult[50][0] ),
  .QN(_05083_)
);

DFF_X1 \sresult[50][10]$_DFFE_PP_  (
  .D(_00610_),
  .CK(clk),
  .Q(\sresult[50][10] ),
  .QN(_05073_)
);

DFF_X1 \sresult[50][11]$_DFFE_PP_  (
  .D(_00611_),
  .CK(clk),
  .Q(\sresult[50][11] ),
  .QN(_05072_)
);

DFF_X1 \sresult[50][1]$_DFFE_PP_  (
  .D(_00601_),
  .CK(clk),
  .Q(\sresult[50][1] ),
  .QN(_05082_)
);

DFF_X1 \sresult[50][2]$_DFFE_PP_  (
  .D(_00602_),
  .CK(clk),
  .Q(\sresult[50][2] ),
  .QN(_05081_)
);

DFF_X1 \sresult[50][3]$_DFFE_PP_  (
  .D(_00603_),
  .CK(clk),
  .Q(\sresult[50][3] ),
  .QN(_05080_)
);

DFF_X1 \sresult[50][4]$_DFFE_PP_  (
  .D(_00604_),
  .CK(clk),
  .Q(\sresult[50][4] ),
  .QN(_05079_)
);

DFF_X1 \sresult[50][5]$_DFFE_PP_  (
  .D(_00605_),
  .CK(clk),
  .Q(\sresult[50][5] ),
  .QN(_05078_)
);

DFF_X1 \sresult[50][6]$_DFFE_PP_  (
  .D(_00606_),
  .CK(clk),
  .Q(\sresult[50][6] ),
  .QN(_05077_)
);

DFF_X1 \sresult[50][7]$_DFFE_PP_  (
  .D(_00607_),
  .CK(clk),
  .Q(\sresult[50][7] ),
  .QN(_05076_)
);

DFF_X1 \sresult[50][8]$_DFFE_PP_  (
  .D(_00608_),
  .CK(clk),
  .Q(\sresult[50][8] ),
  .QN(_05075_)
);

DFF_X1 \sresult[50][9]$_DFFE_PP_  (
  .D(_00609_),
  .CK(clk),
  .Q(\sresult[50][9] ),
  .QN(_05074_)
);

DFF_X1 \sresult[51][0]$_DFFE_PP_  (
  .D(_00612_),
  .CK(clk),
  .Q(\sresult[51][0] ),
  .QN(_05071_)
);

DFF_X1 \sresult[51][10]$_DFFE_PP_  (
  .D(_00622_),
  .CK(clk),
  .Q(\sresult[51][10] ),
  .QN(_05061_)
);

DFF_X1 \sresult[51][11]$_DFFE_PP_  (
  .D(_00623_),
  .CK(clk),
  .Q(\sresult[51][11] ),
  .QN(_05060_)
);

DFF_X1 \sresult[51][1]$_DFFE_PP_  (
  .D(_00613_),
  .CK(clk),
  .Q(\sresult[51][1] ),
  .QN(_05070_)
);

DFF_X1 \sresult[51][2]$_DFFE_PP_  (
  .D(_00614_),
  .CK(clk),
  .Q(\sresult[51][2] ),
  .QN(_05069_)
);

DFF_X1 \sresult[51][3]$_DFFE_PP_  (
  .D(_00615_),
  .CK(clk),
  .Q(\sresult[51][3] ),
  .QN(_05068_)
);

DFF_X1 \sresult[51][4]$_DFFE_PP_  (
  .D(_00616_),
  .CK(clk),
  .Q(\sresult[51][4] ),
  .QN(_05067_)
);

DFF_X1 \sresult[51][5]$_DFFE_PP_  (
  .D(_00617_),
  .CK(clk),
  .Q(\sresult[51][5] ),
  .QN(_05066_)
);

DFF_X1 \sresult[51][6]$_DFFE_PP_  (
  .D(_00618_),
  .CK(clk),
  .Q(\sresult[51][6] ),
  .QN(_05065_)
);

DFF_X1 \sresult[51][7]$_DFFE_PP_  (
  .D(_00619_),
  .CK(clk),
  .Q(\sresult[51][7] ),
  .QN(_05064_)
);

DFF_X1 \sresult[51][8]$_DFFE_PP_  (
  .D(_00620_),
  .CK(clk),
  .Q(\sresult[51][8] ),
  .QN(_05063_)
);

DFF_X1 \sresult[51][9]$_DFFE_PP_  (
  .D(_00621_),
  .CK(clk),
  .Q(\sresult[51][9] ),
  .QN(_05062_)
);

DFF_X1 \sresult[52][0]$_DFFE_PP_  (
  .D(_00624_),
  .CK(clk),
  .Q(\sresult[52][0] ),
  .QN(_05059_)
);

DFF_X1 \sresult[52][10]$_DFFE_PP_  (
  .D(_00634_),
  .CK(clk),
  .Q(\sresult[52][10] ),
  .QN(_05049_)
);

DFF_X1 \sresult[52][11]$_DFFE_PP_  (
  .D(_00635_),
  .CK(clk),
  .Q(\sresult[52][11] ),
  .QN(_05048_)
);

DFF_X1 \sresult[52][1]$_DFFE_PP_  (
  .D(_00625_),
  .CK(clk),
  .Q(\sresult[52][1] ),
  .QN(_05058_)
);

DFF_X1 \sresult[52][2]$_DFFE_PP_  (
  .D(_00626_),
  .CK(clk),
  .Q(\sresult[52][2] ),
  .QN(_05057_)
);

DFF_X1 \sresult[52][3]$_DFFE_PP_  (
  .D(_00627_),
  .CK(clk),
  .Q(\sresult[52][3] ),
  .QN(_05056_)
);

DFF_X1 \sresult[52][4]$_DFFE_PP_  (
  .D(_00628_),
  .CK(clk),
  .Q(\sresult[52][4] ),
  .QN(_05055_)
);

DFF_X1 \sresult[52][5]$_DFFE_PP_  (
  .D(_00629_),
  .CK(clk),
  .Q(\sresult[52][5] ),
  .QN(_05054_)
);

DFF_X1 \sresult[52][6]$_DFFE_PP_  (
  .D(_00630_),
  .CK(clk),
  .Q(\sresult[52][6] ),
  .QN(_05053_)
);

DFF_X1 \sresult[52][7]$_DFFE_PP_  (
  .D(_00631_),
  .CK(clk),
  .Q(\sresult[52][7] ),
  .QN(_05052_)
);

DFF_X1 \sresult[52][8]$_DFFE_PP_  (
  .D(_00632_),
  .CK(clk),
  .Q(\sresult[52][8] ),
  .QN(_05051_)
);

DFF_X1 \sresult[52][9]$_DFFE_PP_  (
  .D(_00633_),
  .CK(clk),
  .Q(\sresult[52][9] ),
  .QN(_05050_)
);

DFF_X1 \sresult[53][0]$_DFFE_PP_  (
  .D(_00636_),
  .CK(clk),
  .Q(\sresult[53][0] ),
  .QN(_05047_)
);

DFF_X1 \sresult[53][10]$_DFFE_PP_  (
  .D(_00646_),
  .CK(clk),
  .Q(\sresult[53][10] ),
  .QN(_05037_)
);

DFF_X1 \sresult[53][11]$_DFFE_PP_  (
  .D(_00647_),
  .CK(clk),
  .Q(\sresult[53][11] ),
  .QN(_05036_)
);

DFF_X1 \sresult[53][1]$_DFFE_PP_  (
  .D(_00637_),
  .CK(clk),
  .Q(\sresult[53][1] ),
  .QN(_05046_)
);

DFF_X1 \sresult[53][2]$_DFFE_PP_  (
  .D(_00638_),
  .CK(clk),
  .Q(\sresult[53][2] ),
  .QN(_05045_)
);

DFF_X1 \sresult[53][3]$_DFFE_PP_  (
  .D(_00639_),
  .CK(clk),
  .Q(\sresult[53][3] ),
  .QN(_05044_)
);

DFF_X1 \sresult[53][4]$_DFFE_PP_  (
  .D(_00640_),
  .CK(clk),
  .Q(\sresult[53][4] ),
  .QN(_05043_)
);

DFF_X1 \sresult[53][5]$_DFFE_PP_  (
  .D(_00641_),
  .CK(clk),
  .Q(\sresult[53][5] ),
  .QN(_05042_)
);

DFF_X1 \sresult[53][6]$_DFFE_PP_  (
  .D(_00642_),
  .CK(clk),
  .Q(\sresult[53][6] ),
  .QN(_05041_)
);

DFF_X1 \sresult[53][7]$_DFFE_PP_  (
  .D(_00643_),
  .CK(clk),
  .Q(\sresult[53][7] ),
  .QN(_05040_)
);

DFF_X1 \sresult[53][8]$_DFFE_PP_  (
  .D(_00644_),
  .CK(clk),
  .Q(\sresult[53][8] ),
  .QN(_05039_)
);

DFF_X1 \sresult[53][9]$_DFFE_PP_  (
  .D(_00645_),
  .CK(clk),
  .Q(\sresult[53][9] ),
  .QN(_05038_)
);

DFF_X1 \sresult[54][0]$_DFFE_PP_  (
  .D(_00648_),
  .CK(clk),
  .Q(\sresult[54][0] ),
  .QN(_05035_)
);

DFF_X1 \sresult[54][10]$_DFFE_PP_  (
  .D(_00658_),
  .CK(clk),
  .Q(\sresult[54][10] ),
  .QN(_05025_)
);

DFF_X1 \sresult[54][11]$_DFFE_PP_  (
  .D(_00659_),
  .CK(clk),
  .Q(\sresult[54][11] ),
  .QN(_05024_)
);

DFF_X1 \sresult[54][1]$_DFFE_PP_  (
  .D(_00649_),
  .CK(clk),
  .Q(\sresult[54][1] ),
  .QN(_05034_)
);

DFF_X1 \sresult[54][2]$_DFFE_PP_  (
  .D(_00650_),
  .CK(clk),
  .Q(\sresult[54][2] ),
  .QN(_05033_)
);

DFF_X1 \sresult[54][3]$_DFFE_PP_  (
  .D(_00651_),
  .CK(clk),
  .Q(\sresult[54][3] ),
  .QN(_05032_)
);

DFF_X1 \sresult[54][4]$_DFFE_PP_  (
  .D(_00652_),
  .CK(clk),
  .Q(\sresult[54][4] ),
  .QN(_05031_)
);

DFF_X1 \sresult[54][5]$_DFFE_PP_  (
  .D(_00653_),
  .CK(clk),
  .Q(\sresult[54][5] ),
  .QN(_05030_)
);

DFF_X1 \sresult[54][6]$_DFFE_PP_  (
  .D(_00654_),
  .CK(clk),
  .Q(\sresult[54][6] ),
  .QN(_05029_)
);

DFF_X1 \sresult[54][7]$_DFFE_PP_  (
  .D(_00655_),
  .CK(clk),
  .Q(\sresult[54][7] ),
  .QN(_05028_)
);

DFF_X1 \sresult[54][8]$_DFFE_PP_  (
  .D(_00656_),
  .CK(clk),
  .Q(\sresult[54][8] ),
  .QN(_05027_)
);

DFF_X1 \sresult[54][9]$_DFFE_PP_  (
  .D(_00657_),
  .CK(clk),
  .Q(\sresult[54][9] ),
  .QN(_05026_)
);

DFF_X1 \sresult[55][0]$_DFFE_PP_  (
  .D(_00660_),
  .CK(clk),
  .Q(\sresult[55][0] ),
  .QN(_05023_)
);

DFF_X1 \sresult[55][10]$_DFFE_PP_  (
  .D(_00670_),
  .CK(clk),
  .Q(\sresult[55][10] ),
  .QN(_05013_)
);

DFF_X1 \sresult[55][11]$_DFFE_PP_  (
  .D(_00671_),
  .CK(clk),
  .Q(\sresult[55][11] ),
  .QN(_05012_)
);

DFF_X1 \sresult[55][1]$_DFFE_PP_  (
  .D(_00661_),
  .CK(clk),
  .Q(\sresult[55][1] ),
  .QN(_05022_)
);

DFF_X1 \sresult[55][2]$_DFFE_PP_  (
  .D(_00662_),
  .CK(clk),
  .Q(\sresult[55][2] ),
  .QN(_05021_)
);

DFF_X1 \sresult[55][3]$_DFFE_PP_  (
  .D(_00663_),
  .CK(clk),
  .Q(\sresult[55][3] ),
  .QN(_05020_)
);

DFF_X1 \sresult[55][4]$_DFFE_PP_  (
  .D(_00664_),
  .CK(clk),
  .Q(\sresult[55][4] ),
  .QN(_05019_)
);

DFF_X1 \sresult[55][5]$_DFFE_PP_  (
  .D(_00665_),
  .CK(clk),
  .Q(\sresult[55][5] ),
  .QN(_05018_)
);

DFF_X1 \sresult[55][6]$_DFFE_PP_  (
  .D(_00666_),
  .CK(clk),
  .Q(\sresult[55][6] ),
  .QN(_05017_)
);

DFF_X1 \sresult[55][7]$_DFFE_PP_  (
  .D(_00667_),
  .CK(clk),
  .Q(\sresult[55][7] ),
  .QN(_05016_)
);

DFF_X1 \sresult[55][8]$_DFFE_PP_  (
  .D(_00668_),
  .CK(clk),
  .Q(\sresult[55][8] ),
  .QN(_05015_)
);

DFF_X1 \sresult[55][9]$_DFFE_PP_  (
  .D(_00669_),
  .CK(clk),
  .Q(\sresult[55][9] ),
  .QN(_05014_)
);

DFF_X1 \sresult[56][0]$_DFFE_PP_  (
  .D(_00672_),
  .CK(clk),
  .Q(\sresult[56][0] ),
  .QN(_05011_)
);

DFF_X1 \sresult[56][10]$_DFFE_PP_  (
  .D(_00682_),
  .CK(clk),
  .Q(\sresult[56][10] ),
  .QN(_05001_)
);

DFF_X1 \sresult[56][11]$_DFFE_PP_  (
  .D(_00683_),
  .CK(clk),
  .Q(\sresult[56][11] ),
  .QN(_05000_)
);

DFF_X1 \sresult[56][1]$_DFFE_PP_  (
  .D(_00673_),
  .CK(clk),
  .Q(\sresult[56][1] ),
  .QN(_05010_)
);

DFF_X1 \sresult[56][2]$_DFFE_PP_  (
  .D(_00674_),
  .CK(clk),
  .Q(\sresult[56][2] ),
  .QN(_05009_)
);

DFF_X1 \sresult[56][3]$_DFFE_PP_  (
  .D(_00675_),
  .CK(clk),
  .Q(\sresult[56][3] ),
  .QN(_05008_)
);

DFF_X1 \sresult[56][4]$_DFFE_PP_  (
  .D(_00676_),
  .CK(clk),
  .Q(\sresult[56][4] ),
  .QN(_05007_)
);

DFF_X1 \sresult[56][5]$_DFFE_PP_  (
  .D(_00677_),
  .CK(clk),
  .Q(\sresult[56][5] ),
  .QN(_05006_)
);

DFF_X1 \sresult[56][6]$_DFFE_PP_  (
  .D(_00678_),
  .CK(clk),
  .Q(\sresult[56][6] ),
  .QN(_05005_)
);

DFF_X1 \sresult[56][7]$_DFFE_PP_  (
  .D(_00679_),
  .CK(clk),
  .Q(\sresult[56][7] ),
  .QN(_05004_)
);

DFF_X1 \sresult[56][8]$_DFFE_PP_  (
  .D(_00680_),
  .CK(clk),
  .Q(\sresult[56][8] ),
  .QN(_05003_)
);

DFF_X1 \sresult[56][9]$_DFFE_PP_  (
  .D(_00681_),
  .CK(clk),
  .Q(\sresult[56][9] ),
  .QN(_05002_)
);

DFF_X1 \sresult[57][0]$_DFFE_PP_  (
  .D(_00684_),
  .CK(clk),
  .Q(\sresult[57][0] ),
  .QN(_04999_)
);

DFF_X1 \sresult[57][10]$_DFFE_PP_  (
  .D(_00694_),
  .CK(clk),
  .Q(\sresult[57][10] ),
  .QN(_04989_)
);

DFF_X1 \sresult[57][11]$_DFFE_PP_  (
  .D(_00695_),
  .CK(clk),
  .Q(\sresult[57][11] ),
  .QN(_04988_)
);

DFF_X1 \sresult[57][1]$_DFFE_PP_  (
  .D(_00685_),
  .CK(clk),
  .Q(\sresult[57][1] ),
  .QN(_04998_)
);

DFF_X1 \sresult[57][2]$_DFFE_PP_  (
  .D(_00686_),
  .CK(clk),
  .Q(\sresult[57][2] ),
  .QN(_04997_)
);

DFF_X1 \sresult[57][3]$_DFFE_PP_  (
  .D(_00687_),
  .CK(clk),
  .Q(\sresult[57][3] ),
  .QN(_04996_)
);

DFF_X1 \sresult[57][4]$_DFFE_PP_  (
  .D(_00688_),
  .CK(clk),
  .Q(\sresult[57][4] ),
  .QN(_04995_)
);

DFF_X1 \sresult[57][5]$_DFFE_PP_  (
  .D(_00689_),
  .CK(clk),
  .Q(\sresult[57][5] ),
  .QN(_04994_)
);

DFF_X1 \sresult[57][6]$_DFFE_PP_  (
  .D(_00690_),
  .CK(clk),
  .Q(\sresult[57][6] ),
  .QN(_04993_)
);

DFF_X1 \sresult[57][7]$_DFFE_PP_  (
  .D(_00691_),
  .CK(clk),
  .Q(\sresult[57][7] ),
  .QN(_04992_)
);

DFF_X1 \sresult[57][8]$_DFFE_PP_  (
  .D(_00692_),
  .CK(clk),
  .Q(\sresult[57][8] ),
  .QN(_04991_)
);

DFF_X1 \sresult[57][9]$_DFFE_PP_  (
  .D(_00693_),
  .CK(clk),
  .Q(\sresult[57][9] ),
  .QN(_04990_)
);

DFF_X1 \sresult[58][0]$_DFFE_PP_  (
  .D(_00696_),
  .CK(clk),
  .Q(\sresult[58][0] ),
  .QN(_04987_)
);

DFF_X1 \sresult[58][10]$_DFFE_PP_  (
  .D(_00706_),
  .CK(clk),
  .Q(\sresult[58][10] ),
  .QN(_04977_)
);

DFF_X1 \sresult[58][11]$_DFFE_PP_  (
  .D(_00707_),
  .CK(clk),
  .Q(\sresult[58][11] ),
  .QN(_04976_)
);

DFF_X1 \sresult[58][1]$_DFFE_PP_  (
  .D(_00697_),
  .CK(clk),
  .Q(\sresult[58][1] ),
  .QN(_04986_)
);

DFF_X1 \sresult[58][2]$_DFFE_PP_  (
  .D(_00698_),
  .CK(clk),
  .Q(\sresult[58][2] ),
  .QN(_04985_)
);

DFF_X1 \sresult[58][3]$_DFFE_PP_  (
  .D(_00699_),
  .CK(clk),
  .Q(\sresult[58][3] ),
  .QN(_04984_)
);

DFF_X1 \sresult[58][4]$_DFFE_PP_  (
  .D(_00700_),
  .CK(clk),
  .Q(\sresult[58][4] ),
  .QN(_04983_)
);

DFF_X1 \sresult[58][5]$_DFFE_PP_  (
  .D(_00701_),
  .CK(clk),
  .Q(\sresult[58][5] ),
  .QN(_04982_)
);

DFF_X1 \sresult[58][6]$_DFFE_PP_  (
  .D(_00702_),
  .CK(clk),
  .Q(\sresult[58][6] ),
  .QN(_04981_)
);

DFF_X1 \sresult[58][7]$_DFFE_PP_  (
  .D(_00703_),
  .CK(clk),
  .Q(\sresult[58][7] ),
  .QN(_04980_)
);

DFF_X1 \sresult[58][8]$_DFFE_PP_  (
  .D(_00704_),
  .CK(clk),
  .Q(\sresult[58][8] ),
  .QN(_04979_)
);

DFF_X1 \sresult[58][9]$_DFFE_PP_  (
  .D(_00705_),
  .CK(clk),
  .Q(\sresult[58][9] ),
  .QN(_04978_)
);

DFF_X1 \sresult[59][0]$_DFFE_PP_  (
  .D(_00708_),
  .CK(clk),
  .Q(\sresult[59][0] ),
  .QN(_04975_)
);

DFF_X1 \sresult[59][10]$_DFFE_PP_  (
  .D(_00718_),
  .CK(clk),
  .Q(\sresult[59][10] ),
  .QN(_04965_)
);

DFF_X1 \sresult[59][11]$_DFFE_PP_  (
  .D(_00719_),
  .CK(clk),
  .Q(\sresult[59][11] ),
  .QN(_04964_)
);

DFF_X1 \sresult[59][1]$_DFFE_PP_  (
  .D(_00709_),
  .CK(clk),
  .Q(\sresult[59][1] ),
  .QN(_04974_)
);

DFF_X1 \sresult[59][2]$_DFFE_PP_  (
  .D(_00710_),
  .CK(clk),
  .Q(\sresult[59][2] ),
  .QN(_04973_)
);

DFF_X1 \sresult[59][3]$_DFFE_PP_  (
  .D(_00711_),
  .CK(clk),
  .Q(\sresult[59][3] ),
  .QN(_04972_)
);

DFF_X1 \sresult[59][4]$_DFFE_PP_  (
  .D(_00712_),
  .CK(clk),
  .Q(\sresult[59][4] ),
  .QN(_04971_)
);

DFF_X1 \sresult[59][5]$_DFFE_PP_  (
  .D(_00713_),
  .CK(clk),
  .Q(\sresult[59][5] ),
  .QN(_04970_)
);

DFF_X1 \sresult[59][6]$_DFFE_PP_  (
  .D(_00714_),
  .CK(clk),
  .Q(\sresult[59][6] ),
  .QN(_04969_)
);

DFF_X1 \sresult[59][7]$_DFFE_PP_  (
  .D(_00715_),
  .CK(clk),
  .Q(\sresult[59][7] ),
  .QN(_04968_)
);

DFF_X1 \sresult[59][8]$_DFFE_PP_  (
  .D(_00716_),
  .CK(clk),
  .Q(\sresult[59][8] ),
  .QN(_04967_)
);

DFF_X1 \sresult[59][9]$_DFFE_PP_  (
  .D(_00717_),
  .CK(clk),
  .Q(\sresult[59][9] ),
  .QN(_04966_)
);

DFF_X1 \sresult[5][0]$_DFFE_PP_  (
  .D(_00060_),
  .CK(clk),
  .Q(\sresult[5][0] ),
  .QN(_05623_)
);

DFF_X1 \sresult[5][10]$_DFFE_PP_  (
  .D(_00070_),
  .CK(clk),
  .Q(\sresult[5][10] ),
  .QN(_05613_)
);

DFF_X1 \sresult[5][11]$_DFFE_PP_  (
  .D(_00071_),
  .CK(clk),
  .Q(\sresult[5][11] ),
  .QN(_05612_)
);

DFF_X1 \sresult[5][1]$_DFFE_PP_  (
  .D(_00061_),
  .CK(clk),
  .Q(\sresult[5][1] ),
  .QN(_05622_)
);

DFF_X1 \sresult[5][2]$_DFFE_PP_  (
  .D(_00062_),
  .CK(clk),
  .Q(\sresult[5][2] ),
  .QN(_05621_)
);

DFF_X1 \sresult[5][3]$_DFFE_PP_  (
  .D(_00063_),
  .CK(clk),
  .Q(\sresult[5][3] ),
  .QN(_05620_)
);

DFF_X1 \sresult[5][4]$_DFFE_PP_  (
  .D(_00064_),
  .CK(clk),
  .Q(\sresult[5][4] ),
  .QN(_05619_)
);

DFF_X1 \sresult[5][5]$_DFFE_PP_  (
  .D(_00065_),
  .CK(clk),
  .Q(\sresult[5][5] ),
  .QN(_05618_)
);

DFF_X1 \sresult[5][6]$_DFFE_PP_  (
  .D(_00066_),
  .CK(clk),
  .Q(\sresult[5][6] ),
  .QN(_05617_)
);

DFF_X1 \sresult[5][7]$_DFFE_PP_  (
  .D(_00067_),
  .CK(clk),
  .Q(\sresult[5][7] ),
  .QN(_05616_)
);

DFF_X1 \sresult[5][8]$_DFFE_PP_  (
  .D(_00068_),
  .CK(clk),
  .Q(\sresult[5][8] ),
  .QN(_05615_)
);

DFF_X1 \sresult[5][9]$_DFFE_PP_  (
  .D(_00069_),
  .CK(clk),
  .Q(\sresult[5][9] ),
  .QN(_05614_)
);

DFF_X1 \sresult[60][0]$_DFFE_PP_  (
  .D(_00720_),
  .CK(clk),
  .Q(\sresult[60][0] ),
  .QN(_04963_)
);

DFF_X1 \sresult[60][10]$_DFFE_PP_  (
  .D(_00730_),
  .CK(clk),
  .Q(\sresult[60][10] ),
  .QN(_04953_)
);

DFF_X1 \sresult[60][11]$_DFFE_PP_  (
  .D(_00731_),
  .CK(clk),
  .Q(\sresult[60][11] ),
  .QN(_04952_)
);

DFF_X1 \sresult[60][1]$_DFFE_PP_  (
  .D(_00721_),
  .CK(clk),
  .Q(\sresult[60][1] ),
  .QN(_04962_)
);

DFF_X1 \sresult[60][2]$_DFFE_PP_  (
  .D(_00722_),
  .CK(clk),
  .Q(\sresult[60][2] ),
  .QN(_04961_)
);

DFF_X1 \sresult[60][3]$_DFFE_PP_  (
  .D(_00723_),
  .CK(clk),
  .Q(\sresult[60][3] ),
  .QN(_04960_)
);

DFF_X1 \sresult[60][4]$_DFFE_PP_  (
  .D(_00724_),
  .CK(clk),
  .Q(\sresult[60][4] ),
  .QN(_04959_)
);

DFF_X1 \sresult[60][5]$_DFFE_PP_  (
  .D(_00725_),
  .CK(clk),
  .Q(\sresult[60][5] ),
  .QN(_04958_)
);

DFF_X1 \sresult[60][6]$_DFFE_PP_  (
  .D(_00726_),
  .CK(clk),
  .Q(\sresult[60][6] ),
  .QN(_04957_)
);

DFF_X1 \sresult[60][7]$_DFFE_PP_  (
  .D(_00727_),
  .CK(clk),
  .Q(\sresult[60][7] ),
  .QN(_04956_)
);

DFF_X1 \sresult[60][8]$_DFFE_PP_  (
  .D(_00728_),
  .CK(clk),
  .Q(\sresult[60][8] ),
  .QN(_04955_)
);

DFF_X1 \sresult[60][9]$_DFFE_PP_  (
  .D(_00729_),
  .CK(clk),
  .Q(\sresult[60][9] ),
  .QN(_04954_)
);

DFF_X1 \sresult[61][0]$_DFFE_PP_  (
  .D(_00732_),
  .CK(clk),
  .Q(\sresult[61][0] ),
  .QN(_04951_)
);

DFF_X1 \sresult[61][10]$_DFFE_PP_  (
  .D(_00742_),
  .CK(clk),
  .Q(\sresult[61][10] ),
  .QN(_04941_)
);

DFF_X1 \sresult[61][11]$_DFFE_PP_  (
  .D(_00743_),
  .CK(clk),
  .Q(\sresult[61][11] ),
  .QN(_04940_)
);

DFF_X1 \sresult[61][1]$_DFFE_PP_  (
  .D(_00733_),
  .CK(clk),
  .Q(\sresult[61][1] ),
  .QN(_04950_)
);

DFF_X1 \sresult[61][2]$_DFFE_PP_  (
  .D(_00734_),
  .CK(clk),
  .Q(\sresult[61][2] ),
  .QN(_04949_)
);

DFF_X1 \sresult[61][3]$_DFFE_PP_  (
  .D(_00735_),
  .CK(clk),
  .Q(\sresult[61][3] ),
  .QN(_04948_)
);

DFF_X1 \sresult[61][4]$_DFFE_PP_  (
  .D(_00736_),
  .CK(clk),
  .Q(\sresult[61][4] ),
  .QN(_04947_)
);

DFF_X1 \sresult[61][5]$_DFFE_PP_  (
  .D(_00737_),
  .CK(clk),
  .Q(\sresult[61][5] ),
  .QN(_04946_)
);

DFF_X1 \sresult[61][6]$_DFFE_PP_  (
  .D(_00738_),
  .CK(clk),
  .Q(\sresult[61][6] ),
  .QN(_04945_)
);

DFF_X1 \sresult[61][7]$_DFFE_PP_  (
  .D(_00739_),
  .CK(clk),
  .Q(\sresult[61][7] ),
  .QN(_04944_)
);

DFF_X1 \sresult[61][8]$_DFFE_PP_  (
  .D(_00740_),
  .CK(clk),
  .Q(\sresult[61][8] ),
  .QN(_04943_)
);

DFF_X1 \sresult[61][9]$_DFFE_PP_  (
  .D(_00741_),
  .CK(clk),
  .Q(\sresult[61][9] ),
  .QN(_04942_)
);

DFF_X1 \sresult[62][0]$_DFFE_PP_  (
  .D(_00744_),
  .CK(clk),
  .Q(\sresult[62][0] ),
  .QN(_04939_)
);

DFF_X1 \sresult[62][10]$_DFFE_PP_  (
  .D(_00754_),
  .CK(clk),
  .Q(\sresult[62][10] ),
  .QN(_04929_)
);

DFF_X1 \sresult[62][11]$_DFFE_PP_  (
  .D(_00755_),
  .CK(clk),
  .Q(\sresult[62][11] ),
  .QN(_04928_)
);

DFF_X1 \sresult[62][1]$_DFFE_PP_  (
  .D(_00745_),
  .CK(clk),
  .Q(\sresult[62][1] ),
  .QN(_04938_)
);

DFF_X1 \sresult[62][2]$_DFFE_PP_  (
  .D(_00746_),
  .CK(clk),
  .Q(\sresult[62][2] ),
  .QN(_04937_)
);

DFF_X1 \sresult[62][3]$_DFFE_PP_  (
  .D(_00747_),
  .CK(clk),
  .Q(\sresult[62][3] ),
  .QN(_04936_)
);

DFF_X1 \sresult[62][4]$_DFFE_PP_  (
  .D(_00748_),
  .CK(clk),
  .Q(\sresult[62][4] ),
  .QN(_04935_)
);

DFF_X1 \sresult[62][5]$_DFFE_PP_  (
  .D(_00749_),
  .CK(clk),
  .Q(\sresult[62][5] ),
  .QN(_04934_)
);

DFF_X1 \sresult[62][6]$_DFFE_PP_  (
  .D(_00750_),
  .CK(clk),
  .Q(\sresult[62][6] ),
  .QN(_04933_)
);

DFF_X1 \sresult[62][7]$_DFFE_PP_  (
  .D(_00751_),
  .CK(clk),
  .Q(\sresult[62][7] ),
  .QN(_04932_)
);

DFF_X1 \sresult[62][8]$_DFFE_PP_  (
  .D(_00752_),
  .CK(clk),
  .Q(\sresult[62][8] ),
  .QN(_04931_)
);

DFF_X1 \sresult[62][9]$_DFFE_PP_  (
  .D(_00753_),
  .CK(clk),
  .Q(\sresult[62][9] ),
  .QN(_04930_)
);

DFF_X1 \sresult[6][0]$_DFFE_PP_  (
  .D(_00072_),
  .CK(clk),
  .Q(\sresult[6][0] ),
  .QN(_05611_)
);

DFF_X1 \sresult[6][10]$_DFFE_PP_  (
  .D(_00082_),
  .CK(clk),
  .Q(\sresult[6][10] ),
  .QN(_05601_)
);

DFF_X1 \sresult[6][11]$_DFFE_PP_  (
  .D(_00083_),
  .CK(clk),
  .Q(\sresult[6][11] ),
  .QN(_05600_)
);

DFF_X1 \sresult[6][1]$_DFFE_PP_  (
  .D(_00073_),
  .CK(clk),
  .Q(\sresult[6][1] ),
  .QN(_05610_)
);

DFF_X1 \sresult[6][2]$_DFFE_PP_  (
  .D(_00074_),
  .CK(clk),
  .Q(\sresult[6][2] ),
  .QN(_05609_)
);

DFF_X1 \sresult[6][3]$_DFFE_PP_  (
  .D(_00075_),
  .CK(clk),
  .Q(\sresult[6][3] ),
  .QN(_05608_)
);

DFF_X1 \sresult[6][4]$_DFFE_PP_  (
  .D(_00076_),
  .CK(clk),
  .Q(\sresult[6][4] ),
  .QN(_05607_)
);

DFF_X1 \sresult[6][5]$_DFFE_PP_  (
  .D(_00077_),
  .CK(clk),
  .Q(\sresult[6][5] ),
  .QN(_05606_)
);

DFF_X1 \sresult[6][6]$_DFFE_PP_  (
  .D(_00078_),
  .CK(clk),
  .Q(\sresult[6][6] ),
  .QN(_05605_)
);

DFF_X1 \sresult[6][7]$_DFFE_PP_  (
  .D(_00079_),
  .CK(clk),
  .Q(\sresult[6][7] ),
  .QN(_05604_)
);

DFF_X1 \sresult[6][8]$_DFFE_PP_  (
  .D(_00080_),
  .CK(clk),
  .Q(\sresult[6][8] ),
  .QN(_05603_)
);

DFF_X1 \sresult[6][9]$_DFFE_PP_  (
  .D(_00081_),
  .CK(clk),
  .Q(\sresult[6][9] ),
  .QN(_05602_)
);

DFF_X1 \sresult[7][0]$_DFFE_PP_  (
  .D(_00084_),
  .CK(clk),
  .Q(\sresult[7][0] ),
  .QN(_05599_)
);

DFF_X1 \sresult[7][10]$_DFFE_PP_  (
  .D(_00094_),
  .CK(clk),
  .Q(\sresult[7][10] ),
  .QN(_05589_)
);

DFF_X1 \sresult[7][11]$_DFFE_PP_  (
  .D(_00095_),
  .CK(clk),
  .Q(\sresult[7][11] ),
  .QN(_05588_)
);

DFF_X1 \sresult[7][1]$_DFFE_PP_  (
  .D(_00085_),
  .CK(clk),
  .Q(\sresult[7][1] ),
  .QN(_05598_)
);

DFF_X1 \sresult[7][2]$_DFFE_PP_  (
  .D(_00086_),
  .CK(clk),
  .Q(\sresult[7][2] ),
  .QN(_05597_)
);

DFF_X1 \sresult[7][3]$_DFFE_PP_  (
  .D(_00087_),
  .CK(clk),
  .Q(\sresult[7][3] ),
  .QN(_05596_)
);

DFF_X1 \sresult[7][4]$_DFFE_PP_  (
  .D(_00088_),
  .CK(clk),
  .Q(\sresult[7][4] ),
  .QN(_05595_)
);

DFF_X1 \sresult[7][5]$_DFFE_PP_  (
  .D(_00089_),
  .CK(clk),
  .Q(\sresult[7][5] ),
  .QN(_05594_)
);

DFF_X1 \sresult[7][6]$_DFFE_PP_  (
  .D(_00090_),
  .CK(clk),
  .Q(\sresult[7][6] ),
  .QN(_05593_)
);

DFF_X1 \sresult[7][7]$_DFFE_PP_  (
  .D(_00091_),
  .CK(clk),
  .Q(\sresult[7][7] ),
  .QN(_05592_)
);

DFF_X1 \sresult[7][8]$_DFFE_PP_  (
  .D(_00092_),
  .CK(clk),
  .Q(\sresult[7][8] ),
  .QN(_05591_)
);

DFF_X1 \sresult[7][9]$_DFFE_PP_  (
  .D(_00093_),
  .CK(clk),
  .Q(\sresult[7][9] ),
  .QN(_05590_)
);

DFF_X1 \sresult[8][0]$_DFFE_PP_  (
  .D(_00096_),
  .CK(clk),
  .Q(\sresult[8][0] ),
  .QN(_05587_)
);

DFF_X1 \sresult[8][10]$_DFFE_PP_  (
  .D(_00106_),
  .CK(clk),
  .Q(\sresult[8][10] ),
  .QN(_05577_)
);

DFF_X1 \sresult[8][11]$_DFFE_PP_  (
  .D(_00107_),
  .CK(clk),
  .Q(\sresult[8][11] ),
  .QN(_05576_)
);

DFF_X1 \sresult[8][1]$_DFFE_PP_  (
  .D(_00097_),
  .CK(clk),
  .Q(\sresult[8][1] ),
  .QN(_05586_)
);

DFF_X1 \sresult[8][2]$_DFFE_PP_  (
  .D(_00098_),
  .CK(clk),
  .Q(\sresult[8][2] ),
  .QN(_05585_)
);

DFF_X1 \sresult[8][3]$_DFFE_PP_  (
  .D(_00099_),
  .CK(clk),
  .Q(\sresult[8][3] ),
  .QN(_05584_)
);

DFF_X1 \sresult[8][4]$_DFFE_PP_  (
  .D(_00100_),
  .CK(clk),
  .Q(\sresult[8][4] ),
  .QN(_05583_)
);

DFF_X1 \sresult[8][5]$_DFFE_PP_  (
  .D(_00101_),
  .CK(clk),
  .Q(\sresult[8][5] ),
  .QN(_05582_)
);

DFF_X1 \sresult[8][6]$_DFFE_PP_  (
  .D(_00102_),
  .CK(clk),
  .Q(\sresult[8][6] ),
  .QN(_05581_)
);

DFF_X1 \sresult[8][7]$_DFFE_PP_  (
  .D(_00103_),
  .CK(clk),
  .Q(\sresult[8][7] ),
  .QN(_05580_)
);

DFF_X1 \sresult[8][8]$_DFFE_PP_  (
  .D(_00104_),
  .CK(clk),
  .Q(\sresult[8][8] ),
  .QN(_05579_)
);

DFF_X1 \sresult[8][9]$_DFFE_PP_  (
  .D(_00105_),
  .CK(clk),
  .Q(\sresult[8][9] ),
  .QN(_05578_)
);

DFF_X1 \sresult[9][0]$_DFFE_PP_  (
  .D(_00108_),
  .CK(clk),
  .Q(\sresult[9][0] ),
  .QN(_05575_)
);

DFF_X1 \sresult[9][10]$_DFFE_PP_  (
  .D(_00118_),
  .CK(clk),
  .Q(\sresult[9][10] ),
  .QN(_05565_)
);

DFF_X1 \sresult[9][11]$_DFFE_PP_  (
  .D(_00119_),
  .CK(clk),
  .Q(\sresult[9][11] ),
  .QN(_05564_)
);

DFF_X1 \sresult[9][1]$_DFFE_PP_  (
  .D(_00109_),
  .CK(clk),
  .Q(\sresult[9][1] ),
  .QN(_05574_)
);

DFF_X1 \sresult[9][2]$_DFFE_PP_  (
  .D(_00110_),
  .CK(clk),
  .Q(\sresult[9][2] ),
  .QN(_05573_)
);

DFF_X1 \sresult[9][3]$_DFFE_PP_  (
  .D(_00111_),
  .CK(clk),
  .Q(\sresult[9][3] ),
  .QN(_05572_)
);

DFF_X1 \sresult[9][4]$_DFFE_PP_  (
  .D(_00112_),
  .CK(clk),
  .Q(\sresult[9][4] ),
  .QN(_05571_)
);

DFF_X1 \sresult[9][5]$_DFFE_PP_  (
  .D(_00113_),
  .CK(clk),
  .Q(\sresult[9][5] ),
  .QN(_05570_)
);

DFF_X1 \sresult[9][6]$_DFFE_PP_  (
  .D(_00114_),
  .CK(clk),
  .Q(\sresult[9][6] ),
  .QN(_05569_)
);

DFF_X1 \sresult[9][7]$_DFFE_PP_  (
  .D(_00115_),
  .CK(clk),
  .Q(\sresult[9][7] ),
  .QN(_05568_)
);

DFF_X1 \sresult[9][8]$_DFFE_PP_  (
  .D(_00116_),
  .CK(clk),
  .Q(\sresult[9][8] ),
  .QN(_05567_)
);

DFF_X1 \sresult[9][9]$_DFFE_PP_  (
  .D(_00117_),
  .CK(clk),
  .Q(\sresult[9][9] ),
  .QN(_05566_)
);
endmodule //zigzag

module jpeg_rzs(input clk, input ena, input rst, input deni, input dci, input [3:0] rleni,
 input [3:0] sizei, input [11:0] ampi, output deno, output dco, output [3:0] rleno, output [3:0] sizeo,
 output [11:0] ampo);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire \amp[0] ;
wire \amp[10] ;
wire \amp[11] ;
wire \amp[1] ;
wire \amp[2] ;
wire \amp[3] ;
wire \amp[4] ;
wire \amp[5] ;
wire \amp[6] ;
wire \amp[7] ;
wire \amp[8] ;
wire \amp[9] ;
wire dc;
wire den;
wire \rlen[0] ;
wire \rlen[1] ;
wire \rlen[2] ;
wire \rlen[3] ;
wire \size[0] ;
wire \size[1] ;
wire \size[2] ;
wire \size[3] ;
wire state;

NAND2_X1 _120_ (
  .A1(rleni[1]),
  .A2(rleni[0]),
  .ZN(_045_)
);

NAND2_X1 _121_ (
  .A1(rleni[3]),
  .A2(rleni[2]),
  .ZN(_046_)
);

NOR2_X1 _122_ (
  .A1(_045_),
  .A2(_046_),
  .ZN(_047_)
);

NOR2_X1 _123_ (
  .A1(sizei[1]),
  .A2(sizei[0]),
  .ZN(_048_)
);

NOR2_X1 _124_ (
  .A1(sizei[3]),
  .A2(sizei[2]),
  .ZN(_049_)
);

NAND3_X1 _125_ (
  .A1(_047_),
  .A2(_048_),
  .A3(_049_),
  .ZN(_050_)
);

BUF_X4 _126_ (
  .A(ena),
  .Z(_051_)
);

NAND2_X4 _127_ (
  .A1(deni),
  .A2(_051_),
  .ZN(_052_)
);

BUF_X8 _128_ (
  .A(_052_),
  .Z(_053_)
);

INV_X1 _129_ (
  .A(_053_),
  .ZN(_054_)
);

NAND2_X1 _130_ (
  .A1(_050_),
  .A2(_054_),
  .ZN(_055_)
);

INV_X1 _131_ (
  .A(state),
  .ZN(_056_)
);

NAND2_X1 _132_ (
  .A1(_056_),
  .A2(_051_),
  .ZN(_057_)
);

NAND3_X1 _133_ (
  .A1(_057_),
  .A2(_053_),
  .A3(den),
  .ZN(_058_)
);

NAND2_X1 _134_ (
  .A1(_055_),
  .A2(_058_),
  .ZN(_000_)
);

NOR2_X1 _135_ (
  .A1(_052_),
  .A2(_056_),
  .ZN(_059_)
);

NOR2_X1 _136_ (
  .A1(rleni[1]),
  .A2(rleni[0]),
  .ZN(_060_)
);

NOR2_X1 _137_ (
  .A1(rleni[3]),
  .A2(rleni[2]),
  .ZN(_061_)
);

INV_X1 _138_ (
  .A(dci),
  .ZN(_062_)
);

NAND3_X1 _139_ (
  .A1(_060_),
  .A2(_061_),
  .A3(_062_),
  .ZN(_063_)
);

NAND2_X1 _140_ (
  .A1(_048_),
  .A2(_049_),
  .ZN(_064_)
);

OAI21_X1 _141_ (
  .A(_059_),
  .B1(_063_),
  .B2(_064_),
  .ZN(_065_)
);

INV_X1 _142_ (
  .A(den),
  .ZN(_066_)
);

INV_X1 _143_ (
  .A(deno),
  .ZN(_067_)
);

OAI22_X1 _144_ (
  .A1(_057_),
  .A2(_066_),
  .B1(_067_),
  .B2(_051_),
  .ZN(_068_)
);

INV_X1 _145_ (
  .A(_068_),
  .ZN(_069_)
);

NAND2_X1 _146_ (
  .A1(_065_),
  .A2(_069_),
  .ZN(_001_)
);

BUF_X4 _147_ (
  .A(_051_),
  .Z(_070_)
);

NOR2_X1 _148_ (
  .A1(_070_),
  .A2(dc),
  .ZN(_071_)
);

AOI21_X1 _149_ (
  .A(_071_),
  .B1(_062_),
  .B2(_070_),
  .ZN(_002_)
);

BUF_X4 _150_ (
  .A(_051_),
  .Z(_072_)
);

MUX2_X1 _151_ (
  .A(rleno[0]),
  .B(\rlen[0] ),
  .S(_072_),
  .Z(_003_)
);

MUX2_X1 _152_ (
  .A(rleno[1]),
  .B(\rlen[1] ),
  .S(_070_),
  .Z(_004_)
);

MUX2_X1 _153_ (
  .A(rleno[2]),
  .B(\rlen[2] ),
  .S(_072_),
  .Z(_005_)
);

MUX2_X1 _154_ (
  .A(rleno[3]),
  .B(\rlen[3] ),
  .S(_070_),
  .Z(_006_)
);

MUX2_X1 _155_ (
  .A(sizeo[0]),
  .B(\size[0] ),
  .S(_072_),
  .Z(_007_)
);

MUX2_X1 _156_ (
  .A(sizeo[1]),
  .B(\size[1] ),
  .S(_051_),
  .Z(_008_)
);

MUX2_X1 _157_ (
  .A(sizeo[2]),
  .B(\size[2] ),
  .S(_051_),
  .Z(_009_)
);

MUX2_X1 _158_ (
  .A(sizeo[3]),
  .B(\size[3] ),
  .S(_070_),
  .Z(_010_)
);

MUX2_X1 _159_ (
  .A(ampo[0]),
  .B(\amp[0] ),
  .S(_072_),
  .Z(_011_)
);

MUX2_X1 _160_ (
  .A(ampo[1]),
  .B(\amp[1] ),
  .S(_072_),
  .Z(_012_)
);

MUX2_X1 _161_ (
  .A(ampo[2]),
  .B(\amp[2] ),
  .S(_070_),
  .Z(_013_)
);

MUX2_X1 _162_ (
  .A(ampo[3]),
  .B(\amp[3] ),
  .S(_072_),
  .Z(_014_)
);

MUX2_X1 _163_ (
  .A(ampo[4]),
  .B(\amp[4] ),
  .S(_070_),
  .Z(_015_)
);

MUX2_X1 _164_ (
  .A(ampo[5]),
  .B(\amp[5] ),
  .S(_072_),
  .Z(_016_)
);

MUX2_X1 _165_ (
  .A(ampo[6]),
  .B(\amp[6] ),
  .S(_070_),
  .Z(_017_)
);

MUX2_X1 _166_ (
  .A(ampo[7]),
  .B(\amp[7] ),
  .S(_072_),
  .Z(_018_)
);

MUX2_X1 _167_ (
  .A(ampo[8]),
  .B(\amp[8] ),
  .S(_072_),
  .Z(_019_)
);

MUX2_X1 _168_ (
  .A(ampo[9]),
  .B(\amp[9] ),
  .S(_070_),
  .Z(_020_)
);

MUX2_X1 _169_ (
  .A(ampo[10]),
  .B(\amp[10] ),
  .S(_072_),
  .Z(_021_)
);

MUX2_X1 _170_ (
  .A(ampo[11]),
  .B(\amp[11] ),
  .S(_070_),
  .Z(_022_)
);

MUX2_X1 _171_ (
  .A(dco),
  .B(dc),
  .S(_051_),
  .Z(_023_)
);

MUX2_X1 _172_ (
  .A(sizei[0]),
  .B(\size[0] ),
  .S(_053_),
  .Z(_024_)
);

BUF_X8 _173_ (
  .A(_052_),
  .Z(_073_)
);

MUX2_X1 _174_ (
  .A(sizei[1]),
  .B(\size[1] ),
  .S(_073_),
  .Z(_025_)
);

MUX2_X1 _175_ (
  .A(sizei[2]),
  .B(\size[2] ),
  .S(_053_),
  .Z(_026_)
);

MUX2_X1 _176_ (
  .A(sizei[3]),
  .B(\size[3] ),
  .S(_053_),
  .Z(_027_)
);

MUX2_X1 _177_ (
  .A(rleni[0]),
  .B(\rlen[0] ),
  .S(_053_),
  .Z(_028_)
);

MUX2_X1 _178_ (
  .A(rleni[1]),
  .B(\rlen[1] ),
  .S(_053_),
  .Z(_029_)
);

MUX2_X1 _179_ (
  .A(rleni[2]),
  .B(\rlen[2] ),
  .S(_053_),
  .Z(_030_)
);

MUX2_X1 _180_ (
  .A(rleni[3]),
  .B(\rlen[3] ),
  .S(_073_),
  .Z(_031_)
);

MUX2_X1 _181_ (
  .A(ampi[0]),
  .B(\amp[0] ),
  .S(_073_),
  .Z(_032_)
);

MUX2_X1 _182_ (
  .A(ampi[1]),
  .B(\amp[1] ),
  .S(_073_),
  .Z(_033_)
);

MUX2_X1 _183_ (
  .A(ampi[2]),
  .B(\amp[2] ),
  .S(_073_),
  .Z(_034_)
);

MUX2_X1 _184_ (
  .A(ampi[3]),
  .B(\amp[3] ),
  .S(_052_),
  .Z(_035_)
);

MUX2_X1 _185_ (
  .A(ampi[4]),
  .B(\amp[4] ),
  .S(_073_),
  .Z(_036_)
);

MUX2_X1 _186_ (
  .A(ampi[5]),
  .B(\amp[5] ),
  .S(_073_),
  .Z(_037_)
);

MUX2_X1 _187_ (
  .A(ampi[6]),
  .B(\amp[6] ),
  .S(_073_),
  .Z(_038_)
);

MUX2_X1 _188_ (
  .A(ampi[7]),
  .B(\amp[7] ),
  .S(_073_),
  .Z(_039_)
);

MUX2_X1 _189_ (
  .A(ampi[8]),
  .B(\amp[8] ),
  .S(_073_),
  .Z(_040_)
);

MUX2_X1 _190_ (
  .A(ampi[9]),
  .B(\amp[9] ),
  .S(_052_),
  .Z(_041_)
);

MUX2_X1 _191_ (
  .A(ampi[10]),
  .B(\amp[10] ),
  .S(_052_),
  .Z(_042_)
);

MUX2_X1 _192_ (
  .A(ampi[11]),
  .B(\amp[11] ),
  .S(_052_),
  .Z(_043_)
);

NAND2_X1 _193_ (
  .A1(_053_),
  .A2(state),
  .ZN(_074_)
);

OAI21_X1 _194_ (
  .A(_074_),
  .B1(_050_),
  .B2(_053_),
  .ZN(_044_)
);

DFF_X1 \amp[0]$_DFFE_PP_  (
  .D(_032_),
  .CK(clk),
  .Q(\amp[0] ),
  .QN(_087_)
);

DFF_X1 \amp[10]$_DFFE_PP_  (
  .D(_042_),
  .CK(clk),
  .Q(\amp[10] ),
  .QN(_077_)
);

DFF_X1 \amp[11]$_DFFE_PP_  (
  .D(_043_),
  .CK(clk),
  .Q(\amp[11] ),
  .QN(_076_)
);

DFF_X1 \amp[1]$_DFFE_PP_  (
  .D(_033_),
  .CK(clk),
  .Q(\amp[1] ),
  .QN(_086_)
);

DFF_X1 \amp[2]$_DFFE_PP_  (
  .D(_034_),
  .CK(clk),
  .Q(\amp[2] ),
  .QN(_085_)
);

DFF_X1 \amp[3]$_DFFE_PP_  (
  .D(_035_),
  .CK(clk),
  .Q(\amp[3] ),
  .QN(_084_)
);

DFF_X1 \amp[4]$_DFFE_PP_  (
  .D(_036_),
  .CK(clk),
  .Q(\amp[4] ),
  .QN(_083_)
);

DFF_X1 \amp[5]$_DFFE_PP_  (
  .D(_037_),
  .CK(clk),
  .Q(\amp[5] ),
  .QN(_082_)
);

DFF_X1 \amp[6]$_DFFE_PP_  (
  .D(_038_),
  .CK(clk),
  .Q(\amp[6] ),
  .QN(_081_)
);

DFF_X1 \amp[7]$_DFFE_PP_  (
  .D(_039_),
  .CK(clk),
  .Q(\amp[7] ),
  .QN(_080_)
);

DFF_X1 \amp[8]$_DFFE_PP_  (
  .D(_040_),
  .CK(clk),
  .Q(\amp[8] ),
  .QN(_079_)
);

DFF_X1 \amp[9]$_DFFE_PP_  (
  .D(_041_),
  .CK(clk),
  .Q(\amp[9] ),
  .QN(_078_)
);

DFF_X1 \ampo[0]$_DFFE_PP_  (
  .D(_011_),
  .CK(clk),
  .Q(ampo[0]),
  .QN(_108_)
);

DFF_X1 \ampo[10]$_DFFE_PP_  (
  .D(_021_),
  .CK(clk),
  .Q(ampo[10]),
  .QN(_098_)
);

DFF_X1 \ampo[11]$_DFFE_PP_  (
  .D(_022_),
  .CK(clk),
  .Q(ampo[11]),
  .QN(_097_)
);

DFF_X1 \ampo[1]$_DFFE_PP_  (
  .D(_012_),
  .CK(clk),
  .Q(ampo[1]),
  .QN(_107_)
);

DFF_X1 \ampo[2]$_DFFE_PP_  (
  .D(_013_),
  .CK(clk),
  .Q(ampo[2]),
  .QN(_106_)
);

DFF_X1 \ampo[3]$_DFFE_PP_  (
  .D(_014_),
  .CK(clk),
  .Q(ampo[3]),
  .QN(_105_)
);

DFF_X1 \ampo[4]$_DFFE_PP_  (
  .D(_015_),
  .CK(clk),
  .Q(ampo[4]),
  .QN(_104_)
);

DFF_X1 \ampo[5]$_DFFE_PP_  (
  .D(_016_),
  .CK(clk),
  .Q(ampo[5]),
  .QN(_103_)
);

DFF_X1 \ampo[6]$_DFFE_PP_  (
  .D(_017_),
  .CK(clk),
  .Q(ampo[6]),
  .QN(_102_)
);

DFF_X1 \ampo[7]$_DFFE_PP_  (
  .D(_018_),
  .CK(clk),
  .Q(ampo[7]),
  .QN(_101_)
);

DFF_X1 \ampo[8]$_DFFE_PP_  (
  .D(_019_),
  .CK(clk),
  .Q(ampo[8]),
  .QN(_100_)
);

DFF_X1 \ampo[9]$_DFFE_PP_  (
  .D(_020_),
  .CK(clk),
  .Q(ampo[9]),
  .QN(_099_)
);

DFF_X1 dc$_DFFE_PP_ (
  .D(_002_),
  .CK(clk),
  .Q(dc),
  .QN(_117_)
);

DFF_X1 dco$_DFFE_PP_ (
  .D(_023_),
  .CK(clk),
  .Q(dco),
  .QN(_096_)
);

DFFR_X1 den$_DFFE_PN0P_ (
  .D(_000_),
  .RN(rst),
  .CK(clk),
  .Q(den),
  .QN(_119_)
);

DFFR_X1 deno$_DFFE_PN0P_ (
  .D(_001_),
  .RN(rst),
  .CK(clk),
  .Q(deno),
  .QN(_118_)
);

DFF_X1 \rlen[0]$_DFFE_PP_  (
  .D(_028_),
  .CK(clk),
  .Q(\rlen[0] ),
  .QN(_091_)
);

DFF_X1 \rlen[1]$_DFFE_PP_  (
  .D(_029_),
  .CK(clk),
  .Q(\rlen[1] ),
  .QN(_090_)
);

DFF_X1 \rlen[2]$_DFFE_PP_  (
  .D(_030_),
  .CK(clk),
  .Q(\rlen[2] ),
  .QN(_089_)
);

DFF_X1 \rlen[3]$_DFFE_PP_  (
  .D(_031_),
  .CK(clk),
  .Q(\rlen[3] ),
  .QN(_088_)
);

DFF_X1 \rleno[0]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(rleno[0]),
  .QN(_116_)
);

DFF_X1 \rleno[1]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(rleno[1]),
  .QN(_115_)
);

DFF_X1 \rleno[2]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(rleno[2]),
  .QN(_114_)
);

DFF_X1 \rleno[3]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(rleno[3]),
  .QN(_113_)
);

DFF_X1 \size[0]$_DFFE_PP_  (
  .D(_024_),
  .CK(clk),
  .Q(\size[0] ),
  .QN(_095_)
);

DFF_X1 \size[1]$_DFFE_PP_  (
  .D(_025_),
  .CK(clk),
  .Q(\size[1] ),
  .QN(_094_)
);

DFF_X1 \size[2]$_DFFE_PP_  (
  .D(_026_),
  .CK(clk),
  .Q(\size[2] ),
  .QN(_093_)
);

DFF_X1 \size[3]$_DFFE_PP_  (
  .D(_027_),
  .CK(clk),
  .Q(\size[3] ),
  .QN(_092_)
);

DFF_X1 \sizeo[0]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(sizeo[0]),
  .QN(_112_)
);

DFF_X1 \sizeo[1]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(sizeo[1]),
  .QN(_111_)
);

DFF_X1 \sizeo[2]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(sizeo[2]),
  .QN(_110_)
);

DFF_X1 \sizeo[3]$_DFFE_PP_  (
  .D(_010_),
  .CK(clk),
  .Q(sizeo[3]),
  .QN(_109_)
);

DFFR_X1 state$_DFFE_PN0P_ (
  .D(_044_),
  .RN(rst),
  .CK(clk),
  .Q(state),
  .QN(_075_)
);
endmodule //jpeg_rzs

module jpeg_rle1(input clk, input rst, input ena, input go, input [11:0] din, output [3:0] rlen,
 output [3:0] size, output [11:0] amp, output den, output dcterm);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire \sample_cnt[0] ;
wire \sample_cnt[1] ;
wire \sample_cnt[2] ;
wire \sample_cnt[3] ;
wire \sample_cnt[4] ;
wire \sample_cnt[5] ;
wire state;
wire \zero_cnt[0] ;
wire \zero_cnt[1] ;
wire \zero_cnt[2] ;
wire \zero_cnt[3] ;

INV_X2 _314_ (
  .A(din[0]),
  .ZN(_305_)
);

INV_X1 _315_ (
  .A(din[1]),
  .ZN(_306_)
);

BUF_X2 _316_ (
  .A(ena),
  .Z(_273_)
);

BUF_X1 _317_ (
  .A(_273_),
  .Z(_274_)
);

NOR2_X1 _318_ (
  .A1(amp[0]),
  .A2(_274_),
  .ZN(_275_)
);

BUF_X2 _319_ (
  .A(din[11]),
  .Z(_276_)
);

BUF_X2 _320_ (
  .A(_276_),
  .Z(_277_)
);

XNOR2_X1 _321_ (
  .A(_277_),
  .B(din[0]),
  .ZN(_039_)
);

BUF_X1 _322_ (
  .A(_273_),
  .Z(_040_)
);

AOI21_X1 _323_ (
  .A(_275_),
  .B1(_039_),
  .B2(_040_),
  .ZN(_007_)
);

INV_X1 _324_ (
  .A(din[11]),
  .ZN(_041_)
);

OR2_X1 _325_ (
  .A1(_041_),
  .A2(_308_),
  .ZN(_042_)
);

OAI21_X1 _326_ (
  .A(_042_),
  .B1(_277_),
  .B2(_306_),
  .ZN(_043_)
);

MUX2_X1 _327_ (
  .A(amp[1]),
  .B(_043_),
  .S(_273_),
  .Z(_008_)
);

INV_X1 _328_ (
  .A(_309_),
  .ZN(_044_)
);

BUF_X4 _329_ (
  .A(din[2]),
  .Z(_045_)
);

NOR2_X2 _330_ (
  .A1(_044_),
  .A2(_045_),
  .ZN(_046_)
);

INV_X1 _331_ (
  .A(_046_),
  .ZN(_047_)
);

NAND2_X1 _332_ (
  .A1(_044_),
  .A2(_045_),
  .ZN(_048_)
);

NAND3_X1 _333_ (
  .A1(_047_),
  .A2(_276_),
  .A3(_048_),
  .ZN(_049_)
);

INV_X2 _334_ (
  .A(_273_),
  .ZN(_050_)
);

BUF_X1 _335_ (
  .A(_041_),
  .Z(_051_)
);

INV_X2 _336_ (
  .A(_045_),
  .ZN(_052_)
);

AOI21_X1 _337_ (
  .A(_050_),
  .B1(_051_),
  .B2(_052_),
  .ZN(_053_)
);

NAND2_X1 _338_ (
  .A1(_049_),
  .A2(_053_),
  .ZN(_054_)
);

INV_X1 _339_ (
  .A(amp[2]),
  .ZN(_055_)
);

OAI21_X1 _340_ (
  .A(_054_),
  .B1(_040_),
  .B2(_055_),
  .ZN(_009_)
);

NOR2_X4 _341_ (
  .A1(_045_),
  .A2(din[1]),
  .ZN(_056_)
);

NAND2_X2 _342_ (
  .A1(_056_),
  .A2(_305_),
  .ZN(_057_)
);

NAND2_X1 _343_ (
  .A1(_057_),
  .A2(din[3]),
  .ZN(_058_)
);

INV_X2 _344_ (
  .A(din[3]),
  .ZN(_059_)
);

NAND3_X1 _345_ (
  .A1(_056_),
  .A2(_059_),
  .A3(_305_),
  .ZN(_060_)
);

NAND3_X1 _346_ (
  .A1(_058_),
  .A2(_060_),
  .A3(_276_),
  .ZN(_061_)
);

AOI21_X1 _347_ (
  .A(_050_),
  .B1(_051_),
  .B2(_059_),
  .ZN(_062_)
);

NAND2_X1 _348_ (
  .A1(_061_),
  .A2(_062_),
  .ZN(_063_)
);

INV_X1 _349_ (
  .A(amp[3]),
  .ZN(_064_)
);

OAI21_X1 _350_ (
  .A(_063_),
  .B1(_040_),
  .B2(_064_),
  .ZN(_010_)
);

BUF_X4 _351_ (
  .A(din[4]),
  .Z(_065_)
);

NOR2_X4 _352_ (
  .A1(din[3]),
  .A2(_065_),
  .ZN(_066_)
);

AOI21_X1 _353_ (
  .A(_041_),
  .B1(_046_),
  .B2(_066_),
  .ZN(_067_)
);

NAND3_X2 _354_ (
  .A1(_052_),
  .A2(_059_),
  .A3(_309_),
  .ZN(_068_)
);

NAND2_X1 _355_ (
  .A1(_068_),
  .A2(_065_),
  .ZN(_069_)
);

AOI21_X1 _356_ (
  .A(_050_),
  .B1(_067_),
  .B2(_069_),
  .ZN(_070_)
);

OAI21_X1 _357_ (
  .A(_070_),
  .B1(_065_),
  .B2(_277_),
  .ZN(_071_)
);

INV_X1 _358_ (
  .A(amp[4]),
  .ZN(_072_)
);

OAI21_X1 _359_ (
  .A(_071_),
  .B1(_040_),
  .B2(_072_),
  .ZN(_011_)
);

NAND4_X1 _360_ (
  .A1(_056_),
  .A2(_066_),
  .A3(din[5]),
  .A4(_305_),
  .ZN(_073_)
);

NAND3_X1 _361_ (
  .A1(_056_),
  .A2(_066_),
  .A3(_305_),
  .ZN(_074_)
);

INV_X1 _362_ (
  .A(din[5]),
  .ZN(_075_)
);

NAND2_X2 _363_ (
  .A1(_074_),
  .A2(_075_),
  .ZN(_076_)
);

NAND2_X1 _364_ (
  .A1(_073_),
  .A2(_076_),
  .ZN(_077_)
);

NAND2_X1 _365_ (
  .A1(_077_),
  .A2(_277_),
  .ZN(_078_)
);

NAND2_X1 _366_ (
  .A1(_075_),
  .A2(_051_),
  .ZN(_079_)
);

NAND3_X1 _367_ (
  .A1(_078_),
  .A2(_274_),
  .A3(_079_),
  .ZN(_080_)
);

INV_X1 _368_ (
  .A(amp[5]),
  .ZN(_081_)
);

OAI21_X1 _369_ (
  .A(_080_),
  .B1(_040_),
  .B2(_081_),
  .ZN(_012_)
);

NOR2_X2 _370_ (
  .A1(din[5]),
  .A2(din[6]),
  .ZN(_082_)
);

NAND3_X1 _371_ (
  .A1(_046_),
  .A2(_066_),
  .A3(_082_),
  .ZN(_083_)
);

NAND2_X1 _372_ (
  .A1(_083_),
  .A2(din[11]),
  .ZN(_084_)
);

INV_X1 _373_ (
  .A(_084_),
  .ZN(_085_)
);

NAND3_X1 _374_ (
  .A1(_046_),
  .A2(_066_),
  .A3(_075_),
  .ZN(_086_)
);

NAND2_X1 _375_ (
  .A1(_086_),
  .A2(din[6]),
  .ZN(_087_)
);

NAND2_X1 _376_ (
  .A1(_085_),
  .A2(_087_),
  .ZN(_088_)
);

INV_X1 _377_ (
  .A(din[6]),
  .ZN(_089_)
);

AOI21_X1 _378_ (
  .A(_050_),
  .B1(_051_),
  .B2(_089_),
  .ZN(_090_)
);

NAND2_X1 _379_ (
  .A1(_088_),
  .A2(_090_),
  .ZN(_091_)
);

INV_X1 _380_ (
  .A(amp[6]),
  .ZN(_092_)
);

OAI21_X1 _381_ (
  .A(_091_),
  .B1(_040_),
  .B2(_092_),
  .ZN(_013_)
);

INV_X1 _382_ (
  .A(din[7]),
  .ZN(_093_)
);

NAND2_X4 _383_ (
  .A1(_066_),
  .A2(_082_),
  .ZN(_094_)
);

OAI21_X2 _384_ (
  .A(_093_),
  .B1(_094_),
  .B2(_057_),
  .ZN(_095_)
);

NOR2_X4 _385_ (
  .A1(_094_),
  .A2(_057_),
  .ZN(_096_)
);

NAND2_X1 _386_ (
  .A1(_096_),
  .A2(din[7]),
  .ZN(_097_)
);

NAND2_X1 _387_ (
  .A1(_095_),
  .A2(_097_),
  .ZN(_098_)
);

NAND2_X1 _388_ (
  .A1(_098_),
  .A2(_277_),
  .ZN(_099_)
);

NAND2_X1 _389_ (
  .A1(_093_),
  .A2(_051_),
  .ZN(_100_)
);

NAND3_X1 _390_ (
  .A1(_099_),
  .A2(_274_),
  .A3(_100_),
  .ZN(_101_)
);

INV_X1 _391_ (
  .A(amp[7]),
  .ZN(_102_)
);

OAI21_X1 _392_ (
  .A(_101_),
  .B1(_040_),
  .B2(_102_),
  .ZN(_014_)
);

NOR2_X1 _393_ (
  .A1(din[5]),
  .A2(_065_),
  .ZN(_103_)
);

NOR2_X1 _394_ (
  .A1(din[7]),
  .A2(din[6]),
  .ZN(_104_)
);

NAND2_X1 _395_ (
  .A1(_103_),
  .A2(_104_),
  .ZN(_105_)
);

NOR2_X2 _396_ (
  .A1(_105_),
  .A2(_068_),
  .ZN(_106_)
);

INV_X1 _397_ (
  .A(din[8]),
  .ZN(_107_)
);

XNOR2_X1 _398_ (
  .A(_106_),
  .B(_107_),
  .ZN(_108_)
);

NAND2_X2 _399_ (
  .A1(_108_),
  .A2(_277_),
  .ZN(_109_)
);

OAI21_X1 _400_ (
  .A(_109_),
  .B1(_107_),
  .B2(_277_),
  .ZN(_110_)
);

MUX2_X1 _401_ (
  .A(amp[8]),
  .B(_110_),
  .S(_274_),
  .Z(_015_)
);

NOR2_X1 _402_ (
  .A1(din[7]),
  .A2(din[8]),
  .ZN(_111_)
);

NAND2_X2 _403_ (
  .A1(_096_),
  .A2(_111_),
  .ZN(_112_)
);

INV_X1 _404_ (
  .A(din[9]),
  .ZN(_113_)
);

NAND2_X2 _405_ (
  .A1(_112_),
  .A2(_113_),
  .ZN(_114_)
);

NAND3_X1 _406_ (
  .A1(_096_),
  .A2(din[9]),
  .A3(_111_),
  .ZN(_115_)
);

NAND3_X2 _407_ (
  .A1(_114_),
  .A2(_115_),
  .A3(_276_),
  .ZN(_116_)
);

OAI21_X1 _408_ (
  .A(_116_),
  .B1(_113_),
  .B2(_277_),
  .ZN(_117_)
);

MUX2_X1 _409_ (
  .A(amp[9]),
  .B(_117_),
  .S(_274_),
  .Z(_016_)
);

INV_X1 _410_ (
  .A(_106_),
  .ZN(_118_)
);

NOR2_X1 _411_ (
  .A1(din[9]),
  .A2(din[8]),
  .ZN(_119_)
);

INV_X1 _412_ (
  .A(_119_),
  .ZN(_120_)
);

OAI21_X1 _413_ (
  .A(din[10]),
  .B1(_118_),
  .B2(_120_),
  .ZN(_121_)
);

INV_X1 _414_ (
  .A(din[10]),
  .ZN(_122_)
);

NAND3_X1 _415_ (
  .A1(_106_),
  .A2(_122_),
  .A3(_119_),
  .ZN(_123_)
);

NAND3_X1 _416_ (
  .A1(_121_),
  .A2(_123_),
  .A3(_277_),
  .ZN(_124_)
);

NAND2_X1 _417_ (
  .A1(_051_),
  .A2(_122_),
  .ZN(_125_)
);

NAND3_X1 _418_ (
  .A1(_124_),
  .A2(_274_),
  .A3(_125_),
  .ZN(_126_)
);

INV_X1 _419_ (
  .A(amp[10]),
  .ZN(_127_)
);

OAI21_X1 _420_ (
  .A(_126_),
  .B1(_040_),
  .B2(_127_),
  .ZN(_017_)
);

NAND2_X1 _421_ (
  .A1(_113_),
  .A2(_051_),
  .ZN(_128_)
);

NAND2_X4 _422_ (
  .A1(_116_),
  .A2(_128_),
  .ZN(_129_)
);

NAND2_X1 _423_ (
  .A1(_107_),
  .A2(_051_),
  .ZN(_130_)
);

NAND2_X2 _424_ (
  .A1(_109_),
  .A2(_130_),
  .ZN(_131_)
);

NAND2_X4 _425_ (
  .A1(_129_),
  .A2(_131_),
  .ZN(_132_)
);

NAND2_X1 _426_ (
  .A1(_051_),
  .A2(din[10]),
  .ZN(_133_)
);

NAND2_X2 _427_ (
  .A1(_124_),
  .A2(_133_),
  .ZN(_134_)
);

NOR2_X4 _428_ (
  .A1(_132_),
  .A2(_134_),
  .ZN(_135_)
);

NAND3_X2 _429_ (
  .A1(_095_),
  .A2(_097_),
  .A3(_276_),
  .ZN(_136_)
);

NAND2_X4 _430_ (
  .A1(_136_),
  .A2(_100_),
  .ZN(_137_)
);

NOR2_X1 _431_ (
  .A1(_089_),
  .A2(_276_),
  .ZN(_138_)
);

AOI21_X4 _432_ (
  .A(_138_),
  .B1(_085_),
  .B2(_087_),
  .ZN(_139_)
);

NAND2_X4 _433_ (
  .A1(_137_),
  .A2(_139_),
  .ZN(_140_)
);

NAND3_X2 _434_ (
  .A1(_073_),
  .A2(_076_),
  .A3(_276_),
  .ZN(_141_)
);

NAND2_X2 _435_ (
  .A1(_141_),
  .A2(_079_),
  .ZN(_142_)
);

INV_X1 _436_ (
  .A(_065_),
  .ZN(_143_)
);

NOR2_X1 _437_ (
  .A1(_143_),
  .A2(_276_),
  .ZN(_144_)
);

AOI21_X2 _438_ (
  .A(_144_),
  .B1(_067_),
  .B2(_069_),
  .ZN(_145_)
);

NAND2_X2 _439_ (
  .A1(_142_),
  .A2(_145_),
  .ZN(_146_)
);

NOR2_X2 _440_ (
  .A1(_140_),
  .A2(_146_),
  .ZN(_147_)
);

NOR2_X1 _441_ (
  .A1(_059_),
  .A2(_276_),
  .ZN(_148_)
);

INV_X1 _442_ (
  .A(_148_),
  .ZN(_149_)
);

NAND2_X1 _443_ (
  .A1(_061_),
  .A2(_149_),
  .ZN(_150_)
);

INV_X1 _444_ (
  .A(_150_),
  .ZN(_151_)
);

OAI21_X1 _445_ (
  .A(_042_),
  .B1(_276_),
  .B2(din[1]),
  .ZN(_152_)
);

NAND2_X1 _446_ (
  .A1(_152_),
  .A2(din[0]),
  .ZN(_153_)
);

NAND2_X1 _447_ (
  .A1(_051_),
  .A2(_045_),
  .ZN(_154_)
);

NAND2_X1 _448_ (
  .A1(_049_),
  .A2(_154_),
  .ZN(_155_)
);

NOR2_X1 _449_ (
  .A1(_153_),
  .A2(_155_),
  .ZN(_156_)
);

INV_X1 _450_ (
  .A(_155_),
  .ZN(_157_)
);

NAND2_X1 _451_ (
  .A1(_157_),
  .A2(_152_),
  .ZN(_158_)
);

OAI21_X1 _452_ (
  .A(_151_),
  .B1(_156_),
  .B2(_158_),
  .ZN(_159_)
);

NAND2_X1 _453_ (
  .A1(_151_),
  .A2(_307_),
  .ZN(_160_)
);

NAND2_X1 _454_ (
  .A1(_159_),
  .A2(_160_),
  .ZN(_161_)
);

NAND3_X2 _455_ (
  .A1(_135_),
  .A2(_147_),
  .A3(_161_),
  .ZN(_162_)
);

NAND2_X1 _456_ (
  .A1(_150_),
  .A2(_145_),
  .ZN(_163_)
);

NAND3_X1 _457_ (
  .A1(_142_),
  .A2(_163_),
  .A3(_139_),
  .ZN(_164_)
);

NAND2_X1 _458_ (
  .A1(_164_),
  .A2(_137_),
  .ZN(_165_)
);

INV_X1 _459_ (
  .A(_140_),
  .ZN(_166_)
);

INV_X1 _460_ (
  .A(_142_),
  .ZN(_167_)
);

NOR2_X1 _461_ (
  .A1(_167_),
  .A2(_145_),
  .ZN(_168_)
);

NAND2_X1 _462_ (
  .A1(_166_),
  .A2(_168_),
  .ZN(_169_)
);

NAND2_X1 _463_ (
  .A1(_165_),
  .A2(_169_),
  .ZN(_170_)
);

NAND2_X2 _464_ (
  .A1(_170_),
  .A2(_135_),
  .ZN(_171_)
);

INV_X1 _465_ (
  .A(_134_),
  .ZN(_172_)
);

NAND2_X1 _466_ (
  .A1(_131_),
  .A2(_137_),
  .ZN(_173_)
);

INV_X1 _467_ (
  .A(_129_),
  .ZN(_174_)
);

OAI21_X1 _468_ (
  .A(_172_),
  .B1(_173_),
  .B2(_174_),
  .ZN(_175_)
);

NAND3_X2 _469_ (
  .A1(_162_),
  .A2(_171_),
  .A3(_175_),
  .ZN(_176_)
);

NAND3_X1 _470_ (
  .A1(_137_),
  .A2(_139_),
  .A3(_142_),
  .ZN(_177_)
);

NAND2_X1 _471_ (
  .A1(_145_),
  .A2(_157_),
  .ZN(_178_)
);

NAND2_X1 _472_ (
  .A1(_163_),
  .A2(_178_),
  .ZN(_179_)
);

NOR2_X1 _473_ (
  .A1(_177_),
  .A2(_179_),
  .ZN(_180_)
);

NAND2_X1 _474_ (
  .A1(_135_),
  .A2(_180_),
  .ZN(_181_)
);

NOR2_X1 _475_ (
  .A1(_134_),
  .A2(_174_),
  .ZN(_182_)
);

INV_X1 _476_ (
  .A(_137_),
  .ZN(_183_)
);

OAI21_X1 _477_ (
  .A(_131_),
  .B1(_183_),
  .B2(_139_),
  .ZN(_184_)
);

NAND2_X1 _478_ (
  .A1(_182_),
  .A2(_184_),
  .ZN(_185_)
);

NAND2_X1 _479_ (
  .A1(_181_),
  .A2(_185_),
  .ZN(_186_)
);

INV_X1 _480_ (
  .A(_135_),
  .ZN(_187_)
);

AND2_X1 _481_ (
  .A1(_151_),
  .A2(_156_),
  .ZN(_188_)
);

NAND2_X1 _482_ (
  .A1(_147_),
  .A2(_188_),
  .ZN(_189_)
);

NOR2_X1 _483_ (
  .A1(_187_),
  .A2(_189_),
  .ZN(_190_)
);

NOR2_X1 _484_ (
  .A1(_186_),
  .A2(_190_),
  .ZN(_191_)
);

NAND2_X1 _485_ (
  .A1(_176_),
  .A2(_191_),
  .ZN(_192_)
);

NOR2_X1 _486_ (
  .A1(_123_),
  .A2(_277_),
  .ZN(_193_)
);

INV_X1 _487_ (
  .A(_193_),
  .ZN(_194_)
);

INV_X1 _488_ (
  .A(state),
  .ZN(_195_)
);

OAI21_X1 _489_ (
  .A(_273_),
  .B1(_194_),
  .B2(_195_),
  .ZN(_196_)
);

INV_X1 _490_ (
  .A(_196_),
  .ZN(_197_)
);

NAND2_X1 _491_ (
  .A1(_192_),
  .A2(_197_),
  .ZN(_198_)
);

BUF_X1 _492_ (
  .A(_050_),
  .Z(_199_)
);

NAND2_X1 _493_ (
  .A1(_199_),
  .A2(size[0]),
  .ZN(_200_)
);

NAND2_X1 _494_ (
  .A1(_198_),
  .A2(_200_),
  .ZN(_018_)
);

AND2_X1 _495_ (
  .A1(_151_),
  .A2(_158_),
  .ZN(_201_)
);

NAND3_X1 _496_ (
  .A1(_135_),
  .A2(_147_),
  .A3(_201_),
  .ZN(_202_)
);

INV_X1 _497_ (
  .A(_139_),
  .ZN(_203_)
);

NOR2_X1 _498_ (
  .A1(_167_),
  .A2(_203_),
  .ZN(_204_)
);

OAI21_X1 _499_ (
  .A(_129_),
  .B1(_173_),
  .B2(_204_),
  .ZN(_205_)
);

NAND2_X1 _500_ (
  .A1(_205_),
  .A2(_172_),
  .ZN(_206_)
);

NAND2_X1 _501_ (
  .A1(_202_),
  .A2(_206_),
  .ZN(_207_)
);

INV_X1 _502_ (
  .A(_207_),
  .ZN(_208_)
);

NAND2_X1 _503_ (
  .A1(_176_),
  .A2(_208_),
  .ZN(_209_)
);

NAND2_X1 _504_ (
  .A1(_209_),
  .A2(_197_),
  .ZN(_210_)
);

NAND2_X1 _505_ (
  .A1(_199_),
  .A2(size[1]),
  .ZN(_211_)
);

NAND2_X1 _506_ (
  .A1(_210_),
  .A2(_211_),
  .ZN(_019_)
);

NAND2_X1 _507_ (
  .A1(_199_),
  .A2(size[2]),
  .ZN(_212_)
);

OAI21_X1 _508_ (
  .A(_212_),
  .B1(_171_),
  .B2(_199_),
  .ZN(_020_)
);

NAND3_X1 _509_ (
  .A1(_162_),
  .A2(_171_),
  .A3(_197_),
  .ZN(_213_)
);

INV_X1 _510_ (
  .A(size[3]),
  .ZN(_214_)
);

OAI21_X1 _511_ (
  .A(_213_),
  .B1(_040_),
  .B2(_214_),
  .ZN(_021_)
);

NAND2_X1 _512_ (
  .A1(_199_),
  .A2(rlen[0]),
  .ZN(_215_)
);

AND3_X1 _513_ (
  .A1(\sample_cnt[2] ),
  .A2(\sample_cnt[3] ),
  .A3(_311_),
  .ZN(_216_)
);

NAND3_X1 _514_ (
  .A1(_216_),
  .A2(\sample_cnt[5] ),
  .A3(\sample_cnt[4] ),
  .ZN(_217_)
);

AOI21_X1 _515_ (
  .A(_217_),
  .B1(_194_),
  .B2(\zero_cnt[0] ),
  .ZN(_218_)
);

NAND2_X1 _516_ (
  .A1(state),
  .A2(_273_),
  .ZN(_219_)
);

INV_X1 _517_ (
  .A(_219_),
  .ZN(_220_)
);

INV_X1 _518_ (
  .A(_217_),
  .ZN(_221_)
);

INV_X1 _519_ (
  .A(_005_),
  .ZN(_222_)
);

OAI21_X1 _520_ (
  .A(_220_),
  .B1(_221_),
  .B2(_222_),
  .ZN(_223_)
);

OAI21_X1 _521_ (
  .A(_215_),
  .B1(_218_),
  .B2(_223_),
  .ZN(_022_)
);

NAND2_X1 _522_ (
  .A1(_199_),
  .A2(rlen[1]),
  .ZN(_224_)
);

AOI21_X1 _523_ (
  .A(_217_),
  .B1(_194_),
  .B2(\zero_cnt[1] ),
  .ZN(_225_)
);

INV_X1 _524_ (
  .A(_000_),
  .ZN(_226_)
);

OAI21_X1 _525_ (
  .A(_220_),
  .B1(_221_),
  .B2(_226_),
  .ZN(_227_)
);

OAI21_X1 _526_ (
  .A(_224_),
  .B1(_225_),
  .B2(_227_),
  .ZN(_023_)
);

NAND2_X1 _527_ (
  .A1(_199_),
  .A2(rlen[2]),
  .ZN(_228_)
);

AOI21_X1 _528_ (
  .A(_217_),
  .B1(_194_),
  .B2(\zero_cnt[2] ),
  .ZN(_229_)
);

INV_X1 _529_ (
  .A(_001_),
  .ZN(_230_)
);

OAI21_X1 _530_ (
  .A(_220_),
  .B1(_221_),
  .B2(_230_),
  .ZN(_231_)
);

OAI21_X1 _531_ (
  .A(_228_),
  .B1(_229_),
  .B2(_231_),
  .ZN(_024_)
);

NAND2_X1 _532_ (
  .A1(_199_),
  .A2(rlen[3]),
  .ZN(_232_)
);

AOI21_X1 _533_ (
  .A(_217_),
  .B1(_194_),
  .B2(\zero_cnt[3] ),
  .ZN(_233_)
);

INV_X1 _534_ (
  .A(_002_),
  .ZN(_234_)
);

OAI21_X1 _535_ (
  .A(_220_),
  .B1(_221_),
  .B2(_234_),
  .ZN(_235_)
);

OAI21_X1 _536_ (
  .A(_232_),
  .B1(_233_),
  .B2(_235_),
  .ZN(_025_)
);

NAND3_X1 _537_ (
  .A1(\zero_cnt[3] ),
  .A2(\zero_cnt[2] ),
  .A3(_312_),
  .ZN(_236_)
);

NAND2_X1 _538_ (
  .A1(_217_),
  .A2(_236_),
  .ZN(_237_)
);

OAI21_X1 _539_ (
  .A(_220_),
  .B1(_194_),
  .B2(_237_),
  .ZN(_238_)
);

NAND2_X1 _540_ (
  .A1(go),
  .A2(_273_),
  .ZN(_239_)
);

INV_X1 _541_ (
  .A(_239_),
  .ZN(_240_)
);

AOI22_X1 _542_ (
  .A1(_240_),
  .A2(_195_),
  .B1(_050_),
  .B2(den),
  .ZN(_241_)
);

NAND2_X1 _543_ (
  .A1(_238_),
  .A2(_241_),
  .ZN(_026_)
);

NAND2_X1 _544_ (
  .A1(_199_),
  .A2(dcterm),
  .ZN(_242_)
);

OAI21_X1 _545_ (
  .A(_242_),
  .B1(_239_),
  .B2(state),
  .ZN(_027_)
);

NOR3_X1 _546_ (
  .A1(_118_),
  .A2(_120_),
  .A3(_125_),
  .ZN(_243_)
);

NAND3_X1 _547_ (
  .A1(_243_),
  .A2(_005_),
  .A3(_274_),
  .ZN(_244_)
);

INV_X1 _548_ (
  .A(\zero_cnt[0] ),
  .ZN(_245_)
);

OAI21_X1 _549_ (
  .A(_244_),
  .B1(_245_),
  .B2(_274_),
  .ZN(_028_)
);

NAND3_X1 _550_ (
  .A1(_243_),
  .A2(_274_),
  .A3(_006_),
  .ZN(_246_)
);

INV_X1 _551_ (
  .A(\zero_cnt[1] ),
  .ZN(_247_)
);

OAI21_X1 _552_ (
  .A(_246_),
  .B1(_247_),
  .B2(_040_),
  .ZN(_029_)
);

NAND2_X1 _553_ (
  .A1(_194_),
  .A2(_273_),
  .ZN(_248_)
);

INV_X1 _554_ (
  .A(_248_),
  .ZN(_249_)
);

NAND2_X1 _555_ (
  .A1(_312_),
  .A2(_273_),
  .ZN(_250_)
);

INV_X1 _556_ (
  .A(\zero_cnt[2] ),
  .ZN(_251_)
);

XNOR2_X1 _557_ (
  .A(_250_),
  .B(_251_),
  .ZN(_252_)
);

NOR2_X1 _558_ (
  .A1(_249_),
  .A2(_252_),
  .ZN(_030_)
);

NAND4_X1 _559_ (
  .A1(\zero_cnt[1] ),
  .A2(_273_),
  .A3(\zero_cnt[2] ),
  .A4(\zero_cnt[0] ),
  .ZN(_253_)
);

XOR2_X1 _560_ (
  .A(_253_),
  .B(\zero_cnt[3] ),
  .Z(_254_)
);

NOR2_X1 _561_ (
  .A1(_249_),
  .A2(_254_),
  .ZN(_031_)
);

NOR2_X1 _562_ (
  .A1(_050_),
  .A2(go),
  .ZN(_255_)
);

INV_X1 _563_ (
  .A(_003_),
  .ZN(_256_)
);

INV_X1 _564_ (
  .A(\sample_cnt[0] ),
  .ZN(_257_)
);

AOI22_X1 _565_ (
  .A1(_255_),
  .A2(_256_),
  .B1(_199_),
  .B2(_257_),
  .ZN(_032_)
);

NAND2_X1 _566_ (
  .A1(_255_),
  .A2(_004_),
  .ZN(_258_)
);

INV_X1 _567_ (
  .A(\sample_cnt[1] ),
  .ZN(_259_)
);

OAI21_X1 _568_ (
  .A(_258_),
  .B1(_259_),
  .B2(_274_),
  .ZN(_033_)
);

INV_X1 _569_ (
  .A(\sample_cnt[2] ),
  .ZN(_260_)
);

INV_X1 _570_ (
  .A(_311_),
  .ZN(_261_)
);

NOR3_X1 _571_ (
  .A1(_260_),
  .A2(_261_),
  .A3(_050_),
  .ZN(_262_)
);

OAI21_X1 _572_ (
  .A(_260_),
  .B1(_261_),
  .B2(_050_),
  .ZN(_263_)
);

INV_X1 _573_ (
  .A(_263_),
  .ZN(_264_)
);

NOR3_X1 _574_ (
  .A1(_262_),
  .A2(_264_),
  .A3(_240_),
  .ZN(_034_)
);

NOR4_X1 _575_ (
  .A1(_260_),
  .A2(_259_),
  .A3(_050_),
  .A4(_257_),
  .ZN(_265_)
);

AND2_X1 _576_ (
  .A1(_265_),
  .A2(\sample_cnt[3] ),
  .ZN(_266_)
);

NOR2_X1 _577_ (
  .A1(_265_),
  .A2(\sample_cnt[3] ),
  .ZN(_267_)
);

NOR3_X1 _578_ (
  .A1(_266_),
  .A2(_267_),
  .A3(_240_),
  .ZN(_035_)
);

AND3_X1 _579_ (
  .A1(_262_),
  .A2(\sample_cnt[3] ),
  .A3(\sample_cnt[4] ),
  .ZN(_268_)
);

AOI21_X1 _580_ (
  .A(\sample_cnt[4] ),
  .B1(_262_),
  .B2(\sample_cnt[3] ),
  .ZN(_269_)
);

NOR3_X1 _581_ (
  .A1(_268_),
  .A2(_269_),
  .A3(_240_),
  .ZN(_036_)
);

NAND2_X1 _582_ (
  .A1(_266_),
  .A2(\sample_cnt[4] ),
  .ZN(_270_)
);

INV_X1 _583_ (
  .A(_270_),
  .ZN(_271_)
);

OAI21_X1 _584_ (
  .A(_239_),
  .B1(_271_),
  .B2(\sample_cnt[5] ),
  .ZN(_272_)
);

AOI21_X1 _585_ (
  .A(_272_),
  .B1(_271_),
  .B2(\sample_cnt[5] ),
  .ZN(_037_)
);

AOI22_X1 _586_ (
  .A1(_221_),
  .A2(_220_),
  .B1(_195_),
  .B2(_239_),
  .ZN(_038_)
);

HA_X1 _587_ (
  .A(_305_),
  .B(_306_),
  .CO(_307_),
  .S(_308_)
);

HA_X1 _588_ (
  .A(_305_),
  .B(_306_),
  .CO(_309_),
  .S(_310_)
);

HA_X1 _589_ (
  .A(\sample_cnt[0] ),
  .B(\sample_cnt[1] ),
  .CO(_311_),
  .S(_004_)
);

HA_X1 _590_ (
  .A(\zero_cnt[0] ),
  .B(\zero_cnt[1] ),
  .CO(_312_),
  .S(_006_)
);

DFF_X1 \amp[0]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(amp[0]),
  .QN(_304_)
);

DFF_X1 \amp[10]$_DFFE_PP_  (
  .D(_017_),
  .CK(clk),
  .Q(amp[10]),
  .QN(_294_)
);

DFF_X1 \amp[1]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(amp[1]),
  .QN(_303_)
);

DFF_X1 \amp[2]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(amp[2]),
  .QN(_302_)
);

DFF_X1 \amp[3]$_DFFE_PP_  (
  .D(_010_),
  .CK(clk),
  .Q(amp[3]),
  .QN(_301_)
);

DFF_X1 \amp[4]$_DFFE_PP_  (
  .D(_011_),
  .CK(clk),
  .Q(amp[4]),
  .QN(_300_)
);

DFF_X1 \amp[5]$_DFFE_PP_  (
  .D(_012_),
  .CK(clk),
  .Q(amp[5]),
  .QN(_299_)
);

DFF_X1 \amp[6]$_DFFE_PP_  (
  .D(_013_),
  .CK(clk),
  .Q(amp[6]),
  .QN(_298_)
);

DFF_X1 \amp[7]$_DFFE_PP_  (
  .D(_014_),
  .CK(clk),
  .Q(amp[7]),
  .QN(_297_)
);

DFF_X1 \amp[8]$_DFFE_PP_  (
  .D(_015_),
  .CK(clk),
  .Q(amp[8]),
  .QN(_296_)
);

DFF_X1 \amp[9]$_DFFE_PP_  (
  .D(_016_),
  .CK(clk),
  .Q(amp[9]),
  .QN(_295_)
);

DFFR_X1 dcterm$_DFFE_PN0P_ (
  .D(_027_),
  .RN(rst),
  .CK(clk),
  .Q(dcterm),
  .QN(_284_)
);

DFFR_X1 den$_DFFE_PN0P_ (
  .D(_026_),
  .RN(rst),
  .CK(clk),
  .Q(den),
  .QN(_285_)
);

DFFR_X1 \rlen[0]$_DFFE_PN0P_  (
  .D(_022_),
  .RN(rst),
  .CK(clk),
  .Q(rlen[0]),
  .QN(_289_)
);

DFFR_X1 \rlen[1]$_DFFE_PN0P_  (
  .D(_023_),
  .RN(rst),
  .CK(clk),
  .Q(rlen[1]),
  .QN(_288_)
);

DFFR_X1 \rlen[2]$_DFFE_PN0P_  (
  .D(_024_),
  .RN(rst),
  .CK(clk),
  .Q(rlen[2]),
  .QN(_287_)
);

DFFR_X1 \rlen[3]$_DFFE_PN0P_  (
  .D(_025_),
  .RN(rst),
  .CK(clk),
  .Q(rlen[3]),
  .QN(_286_)
);

DFF_X1 \sample_cnt[0]$_SDFFCE_PP1P_  (
  .D(_032_),
  .CK(clk),
  .Q(\sample_cnt[0] ),
  .QN(_003_)
);

DFF_X1 \sample_cnt[1]$_SDFFCE_PP0P_  (
  .D(_033_),
  .CK(clk),
  .Q(\sample_cnt[1] ),
  .QN(_283_)
);

DFF_X1 \sample_cnt[2]$_SDFFCE_PP0P_  (
  .D(_034_),
  .CK(clk),
  .Q(\sample_cnt[2] ),
  .QN(_282_)
);

DFF_X1 \sample_cnt[3]$_SDFFCE_PP0P_  (
  .D(_035_),
  .CK(clk),
  .Q(\sample_cnt[3] ),
  .QN(_281_)
);

DFF_X1 \sample_cnt[4]$_SDFFCE_PP0P_  (
  .D(_036_),
  .CK(clk),
  .Q(\sample_cnt[4] ),
  .QN(_280_)
);

DFF_X1 \sample_cnt[5]$_SDFFCE_PP0P_  (
  .D(_037_),
  .CK(clk),
  .Q(\sample_cnt[5] ),
  .QN(_279_)
);

DFFR_X1 \size[0]$_DFFE_PN0P_  (
  .D(_018_),
  .RN(rst),
  .CK(clk),
  .Q(size[0]),
  .QN(_293_)
);

DFFR_X1 \size[1]$_DFFE_PN0P_  (
  .D(_019_),
  .RN(rst),
  .CK(clk),
  .Q(size[1]),
  .QN(_292_)
);

DFFR_X1 \size[2]$_DFFE_PN0P_  (
  .D(_020_),
  .RN(rst),
  .CK(clk),
  .Q(size[2]),
  .QN(_291_)
);

DFFR_X1 \size[3]$_DFFE_PN0P_  (
  .D(_021_),
  .RN(rst),
  .CK(clk),
  .Q(size[3]),
  .QN(_290_)
);

DFFR_X1 state$_DFFE_PN0P_ (
  .D(_038_),
  .RN(rst),
  .CK(clk),
  .Q(state),
  .QN(_278_)
);

DFF_X1 \zero_cnt[0]$_SDFFCE_PP0P_  (
  .D(_028_),
  .CK(clk),
  .Q(\zero_cnt[0] ),
  .QN(_005_)
);

DFF_X1 \zero_cnt[1]$_SDFFCE_PP0P_  (
  .D(_029_),
  .CK(clk),
  .Q(\zero_cnt[1] ),
  .QN(_000_)
);

DFF_X1 \zero_cnt[2]$_SDFFCE_PP0P_  (
  .D(_030_),
  .CK(clk),
  .Q(\zero_cnt[2] ),
  .QN(_001_)
);

DFF_X1 \zero_cnt[3]$_SDFFCE_PP0P_  (
  .D(_031_),
  .CK(clk),
  .Q(\zero_cnt[3] ),
  .QN(_002_)
);
endmodule //jpeg_rle1

module \$paramod$ee2aa8736952ca7eee7f4751cab786a479da4583\div_uu (input clk, input ena,
 input [23:0] z, input [11:0] d, output [11:0] q, output [11:0] s, output div0, output ovf);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire _0032_;
wire _0033_;
wire _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire _0066_;
wire _0067_;
wire _0068_;
wire _0069_;
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
wire _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
wire _0444_;
wire _0445_;
wire _0446_;
wire _0447_;
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire _0658_;
wire _0659_;
wire _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire _0673_;
wire _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire _0679_;
wire _0680_;
wire _0681_;
wire _0682_;
wire _0683_;
wire _0684_;
wire _0685_;
wire _0686_;
wire _0687_;
wire _0688_;
wire _0689_;
wire _0690_;
wire _0691_;
wire _0692_;
wire _0693_;
wire _0694_;
wire _0695_;
wire _0696_;
wire _0697_;
wire _0698_;
wire _0699_;
wire _0700_;
wire _0701_;
wire _0702_;
wire _0703_;
wire _0704_;
wire _0705_;
wire _0706_;
wire _0707_;
wire _0708_;
wire _0709_;
wire _0710_;
wire _0711_;
wire _0712_;
wire _0713_;
wire _0714_;
wire _0715_;
wire _0716_;
wire _0717_;
wire _0718_;
wire _0719_;
wire _0720_;
wire _0721_;
wire _0722_;
wire _0723_;
wire _0724_;
wire _0725_;
wire _0726_;
wire _0727_;
wire _0728_;
wire _0729_;
wire _0730_;
wire _0731_;
wire _0732_;
wire _0733_;
wire _0734_;
wire _0735_;
wire _0736_;
wire _0737_;
wire _0738_;
wire _0739_;
wire _0740_;
wire _0741_;
wire _0742_;
wire _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0748_;
wire _0749_;
wire _0750_;
wire _0751_;
wire _0752_;
wire _0753_;
wire _0754_;
wire _0755_;
wire _0756_;
wire _0757_;
wire _0758_;
wire _0759_;
wire _0760_;
wire _0761_;
wire _0762_;
wire _0763_;
wire _0764_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire _0780_;
wire _0781_;
wire _0782_;
wire _0783_;
wire _0784_;
wire _0785_;
wire _0786_;
wire _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire _0795_;
wire _0796_;
wire _0797_;
wire _0798_;
wire _0799_;
wire _0800_;
wire _0801_;
wire _0802_;
wire _0803_;
wire _0804_;
wire _0805_;
wire _0806_;
wire _0807_;
wire _0808_;
wire _0809_;
wire _0810_;
wire _0811_;
wire _0812_;
wire _0813_;
wire _0814_;
wire _0815_;
wire _0816_;
wire _0817_;
wire _0818_;
wire _0819_;
wire _0820_;
wire _0821_;
wire _0822_;
wire _0823_;
wire _0824_;
wire _0825_;
wire _0826_;
wire _0827_;
wire _0828_;
wire _0829_;
wire _0830_;
wire _0831_;
wire _0832_;
wire _0833_;
wire _0834_;
wire _0835_;
wire _0836_;
wire _0837_;
wire _0838_;
wire _0839_;
wire _0840_;
wire _0841_;
wire _0842_;
wire _0843_;
wire _0844_;
wire _0845_;
wire _0846_;
wire _0847_;
wire _0848_;
wire _0849_;
wire _0850_;
wire _0851_;
wire _0852_;
wire _0853_;
wire _0854_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0858_;
wire _0859_;
wire _0860_;
wire _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0865_;
wire _0866_;
wire _0867_;
wire _0868_;
wire _0869_;
wire _0870_;
wire _0871_;
wire _0872_;
wire _0873_;
wire _0874_;
wire _0875_;
wire _0876_;
wire _0877_;
wire _0878_;
wire _0879_;
wire _0880_;
wire _0881_;
wire _0882_;
wire _0883_;
wire _0884_;
wire _0885_;
wire _0886_;
wire _0887_;
wire _0888_;
wire _0889_;
wire _0890_;
wire _0891_;
wire _0892_;
wire _0893_;
wire _0894_;
wire _0895_;
wire _0896_;
wire _0897_;
wire _0898_;
wire _0899_;
wire _0900_;
wire _0901_;
wire _0902_;
wire _0903_;
wire _0904_;
wire _0905_;
wire _0906_;
wire _0907_;
wire _0908_;
wire _0909_;
wire _0910_;
wire _0911_;
wire _0912_;
wire _0913_;
wire _0914_;
wire _0915_;
wire _0916_;
wire _0917_;
wire _0918_;
wire _0919_;
wire _0920_;
wire _0921_;
wire _0922_;
wire _0923_;
wire _0924_;
wire _0925_;
wire _0926_;
wire _0927_;
wire _0928_;
wire _0929_;
wire _0930_;
wire _0931_;
wire _0932_;
wire _0933_;
wire _0934_;
wire _0935_;
wire _0936_;
wire _0937_;
wire _0938_;
wire _0939_;
wire _0940_;
wire _0941_;
wire _0942_;
wire _0943_;
wire _0944_;
wire _0945_;
wire _0946_;
wire _0947_;
wire _0948_;
wire _0949_;
wire _0950_;
wire _0951_;
wire _0952_;
wire _0953_;
wire _0954_;
wire _0955_;
wire _0956_;
wire _0957_;
wire _0958_;
wire _0959_;
wire _0960_;
wire _0961_;
wire _0962_;
wire _0963_;
wire _0964_;
wire _0965_;
wire _0966_;
wire _0967_;
wire _0968_;
wire _0969_;
wire _0970_;
wire _0971_;
wire _0972_;
wire _0973_;
wire _0974_;
wire _0975_;
wire _0976_;
wire _0977_;
wire _0978_;
wire _0979_;
wire _0980_;
wire _0981_;
wire _0982_;
wire _0983_;
wire _0984_;
wire _0985_;
wire _0986_;
wire _0987_;
wire _0988_;
wire _0989_;
wire _0990_;
wire _0991_;
wire _0992_;
wire _0993_;
wire _0994_;
wire _0995_;
wire _0996_;
wire _0997_;
wire _0998_;
wire _0999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire _1235_;
wire _1236_;
wire _1237_;
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
wire _1246_;
wire _1247_;
wire _1248_;
wire _1249_;
wire _1250_;
wire _1251_;
wire _1252_;
wire _1253_;
wire _1254_;
wire _1255_;
wire _1256_;
wire _1257_;
wire _1258_;
wire _1259_;
wire _1260_;
wire _1261_;
wire _1262_;
wire _1263_;
wire _1264_;
wire _1265_;
wire _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
wire _1270_;
wire _1271_;
wire _1272_;
wire _1273_;
wire _1274_;
wire _1275_;
wire _1276_;
wire _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire _1283_;
wire _1284_;
wire _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire _1291_;
wire _1292_;
wire _1293_;
wire _1294_;
wire _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1346_;
wire _1347_;
wire _1348_;
wire _1350_;
wire _1351_;
wire _1353_;
wire _1361_;
wire _1363_;
wire _1364_;
wire _1366_;
wire _1367_;
wire _1368_;
wire _1369_;
wire _1371_;
wire _1373_;
wire _1379_;
wire _1381_;
wire _1383_;
wire _1384_;
wire _1385_;
wire _1386_;
wire _1397_;
wire _1404_;
wire _1406_;
wire _1408_;
wire _1410_;
wire _1411_;
wire _1413_;
wire _1414_;
wire _1415_;
wire _1416_;
wire _1417_;
wire _1418_;
wire _1426_;
wire _1427_;
wire _1435_;
wire _1444_;
wire _1446_;
wire _1447_;
wire _1449_;
wire _1455_;
wire _1458_;
wire _1460_;
wire _1461_;
wire _1477_;
wire _1485_;
wire _1490_;
wire _1492_;
wire _1493_;
wire _1494_;
wire _1495_;
wire _1496_;
wire _1497_;
wire _1498_;
wire _1499_;
wire _1500_;
wire _1501_;
wire _1502_;
wire _1503_;
wire _1504_;
wire _1505_;
wire _1506_;
wire _1507_;
wire _1508_;
wire _1509_;
wire _1510_;
wire _1511_;
wire _1512_;
wire _1513_;
wire _1514_;
wire _1515_;
wire _1516_;
wire _1517_;
wire _1518_;
wire _1519_;
wire _1520_;
wire _1521_;
wire _1522_;
wire _1523_;
wire _1524_;
wire _1525_;
wire _1526_;
wire _1527_;
wire _1528_;
wire _1529_;
wire _1530_;
wire _1531_;
wire _1532_;
wire _1533_;
wire _1534_;
wire _1535_;
wire _1536_;
wire _1537_;
wire _1538_;
wire _1539_;
wire _1540_;
wire _1541_;
wire _1542_;
wire _1543_;
wire _1544_;
wire _1545_;
wire _1546_;
wire _1547_;
wire _1548_;
wire _1549_;
wire _1550_;
wire _1551_;
wire _1552_;
wire _1553_;
wire _1554_;
wire _1555_;
wire _1556_;
wire _1557_;
wire _1558_;
wire _1559_;
wire _1560_;
wire _1561_;
wire _1562_;
wire _1563_;
wire _1564_;
wire _1565_;
wire _1566_;
wire _1567_;
wire _1568_;
wire _1569_;
wire _1570_;
wire _1571_;
wire _1572_;
wire _1573_;
wire _1574_;
wire _1575_;
wire _1576_;
wire _1577_;
wire _1578_;
wire _1579_;
wire _1580_;
wire _1581_;
wire _1582_;
wire _1583_;
wire _1584_;
wire _1585_;
wire _1586_;
wire _1587_;
wire _1588_;
wire _1589_;
wire _1590_;
wire _1591_;
wire _1592_;
wire _1593_;
wire _1594_;
wire _1595_;
wire _1596_;
wire _1597_;
wire _1598_;
wire _1599_;
wire _1600_;
wire _1601_;
wire _1602_;
wire _1603_;
wire _1604_;
wire _1605_;
wire _1606_;
wire _1607_;
wire _1608_;
wire _1609_;
wire _1610_;
wire _1611_;
wire _1612_;
wire _1613_;
wire _1614_;
wire _1615_;
wire _1616_;
wire _1617_;
wire _1618_;
wire _1619_;
wire _1620_;
wire _1621_;
wire _1622_;
wire _1623_;
wire _1624_;
wire _1625_;
wire _1626_;
wire _1627_;
wire _1628_;
wire _1629_;
wire _1630_;
wire _1631_;
wire _1632_;
wire _1633_;
wire _1634_;
wire _1635_;
wire _1636_;
wire _1637_;
wire _1638_;
wire _1639_;
wire _1640_;
wire _1641_;
wire _1642_;
wire _1643_;
wire _1644_;
wire _1645_;
wire _1646_;
wire _1647_;
wire _1648_;
wire _1649_;
wire _1650_;
wire _1651_;
wire _1652_;
wire _1653_;
wire _1654_;
wire _1655_;
wire _1656_;
wire _1657_;
wire _1658_;
wire _1659_;
wire _1660_;
wire _1661_;
wire _1662_;
wire _1663_;
wire _1664_;
wire _1665_;
wire _1666_;
wire _1667_;
wire _1668_;
wire _1669_;
wire _1670_;
wire _1671_;
wire _1672_;
wire _1673_;
wire _1674_;
wire _1675_;
wire _1676_;
wire _1677_;
wire _1678_;
wire _1679_;
wire _1680_;
wire _1681_;
wire _1682_;
wire _1683_;
wire _1684_;
wire _1685_;
wire _1686_;
wire _1687_;
wire _1688_;
wire _1689_;
wire _1690_;
wire _1691_;
wire _1692_;
wire _1693_;
wire _1694_;
wire _1695_;
wire _1696_;
wire _1697_;
wire _1698_;
wire _1699_;
wire _1700_;
wire _1701_;
wire _1702_;
wire _1703_;
wire _1704_;
wire _1705_;
wire _1706_;
wire _1707_;
wire _1708_;
wire _1709_;
wire _1710_;
wire _1711_;
wire _1712_;
wire _1713_;
wire _1714_;
wire _1715_;
wire _1716_;
wire _1717_;
wire _1718_;
wire _1719_;
wire _1720_;
wire _1721_;
wire _1722_;
wire _1723_;
wire _1724_;
wire _1725_;
wire _1726_;
wire _1727_;
wire _1728_;
wire _1729_;
wire _1859_;
wire _1861_;
wire _1862_;
wire _1863_;
wire _1864_;
wire _1865_;
wire _1866_;
wire _1867_;
wire _1868_;
wire _1869_;
wire _1870_;
wire _1871_;
wire _1872_;
wire _1873_;
wire _1874_;
wire _1875_;
wire _1876_;
wire _1877_;
wire _1878_;
wire _1879_;
wire _1880_;
wire _1881_;
wire _1882_;
wire _1883_;
wire _1884_;
wire _1885_;
wire _1893_;
wire _1897_;
wire _1898_;
wire _1899_;
wire _1901_;
wire _1933_;
wire _1934_;
wire _1936_;
wire _1937_;
wire _1938_;
wire _1939_;
wire _1940_;
wire _1941_;
wire _1942_;
wire _1943_;
wire _1944_;
wire _1945_;
wire _1946_;
wire _1947_;
wire _1948_;
wire _1949_;
wire _1950_;
wire _1951_;
wire _1952_;
wire _1953_;
wire _1954_;
wire _1955_;
wire _1956_;
wire _1957_;
wire _1958_;
wire _1959_;
wire _1960_;
wire _1961_;
wire _1962_;
wire _1963_;
wire _1964_;
wire _1965_;
wire _1966_;
wire _1967_;
wire _1968_;
wire _1969_;
wire _1970_;
wire _1971_;
wire _1972_;
wire _1973_;
wire _1974_;
wire _1975_;
wire _1976_;
wire _1977_;
wire _1978_;
wire _1979_;
wire _1980_;
wire _1981_;
wire _1982_;
wire _1983_;
wire _1984_;
wire _1985_;
wire _1986_;
wire _1987_;
wire _1988_;
wire _1989_;
wire _1990_;
wire _1991_;
wire _1992_;
wire _1993_;
wire _1994_;
wire _1995_;
wire _1996_;
wire _1997_;
wire _1998_;
wire _1999_;
wire _2000_;
wire _2001_;
wire _2002_;
wire _2003_;
wire _2004_;
wire _2005_;
wire _2006_;
wire _2007_;
wire _2008_;
wire _2009_;
wire _2010_;
wire _2011_;
wire _2012_;
wire _2013_;
wire _2014_;
wire _2015_;
wire _2016_;
wire _2017_;
wire _2018_;
wire _2019_;
wire _2020_;
wire _2021_;
wire _2022_;
wire _2023_;
wire _2024_;
wire _2025_;
wire _2026_;
wire _2027_;
wire _2028_;
wire _2029_;
wire _2030_;
wire _2031_;
wire _2032_;
wire _2033_;
wire _2034_;
wire _2035_;
wire _2036_;
wire _2037_;
wire _2038_;
wire _2039_;
wire _2040_;
wire _2041_;
wire _2042_;
wire _2043_;
wire _2044_;
wire _2045_;
wire _2046_;
wire _2047_;
wire _2048_;
wire _2049_;
wire _2050_;
wire _2051_;
wire _2052_;
wire _2054_;
wire _2057_;
wire _2066_;
wire _2067_;
wire _2068_;
wire _2069_;
wire _2070_;
wire _2071_;
wire _2072_;
wire _2073_;
wire _2074_;
wire _2075_;
wire _2076_;
wire _2077_;
wire _2078_;
wire _2079_;
wire _2080_;
wire _2081_;
wire _2082_;
wire _2083_;
wire _2084_;
wire _2085_;
wire _2086_;
wire _2087_;
wire _2088_;
wire _2089_;
wire _2090_;
wire _2091_;
wire _2092_;
wire _2093_;
wire _2094_;
wire _2095_;
wire _2096_;
wire _2097_;
wire _2098_;
wire _2099_;
wire _2100_;
wire _2101_;
wire _2102_;
wire _2103_;
wire _2104_;
wire _2105_;
wire _2106_;
wire _2107_;
wire _2108_;
wire _2109_;
wire _2110_;
wire _2111_;
wire _2112_;
wire _2113_;
wire _2114_;
wire _2115_;
wire _2116_;
wire _2117_;
wire _2118_;
wire _2119_;
wire _2120_;
wire _2121_;
wire _2122_;
wire _2123_;
wire _2124_;
wire _2125_;
wire _2126_;
wire _2127_;
wire _2128_;
wire _2129_;
wire _2130_;
wire _2131_;
wire _2132_;
wire _2133_;
wire _2134_;
wire _2135_;
wire _2136_;
wire _2137_;
wire _2138_;
wire _2139_;
wire _2140_;
wire _2141_;
wire _2142_;
wire _2143_;
wire _2144_;
wire _2145_;
wire _2146_;
wire _2147_;
wire _2148_;
wire _2149_;
wire _2150_;
wire _2151_;
wire _2152_;
wire _2153_;
wire _2154_;
wire _2155_;
wire _2156_;
wire _2157_;
wire _2158_;
wire _2159_;
wire _2160_;
wire _2161_;
wire _2162_;
wire _2163_;
wire _2164_;
wire _2165_;
wire _2166_;
wire _2167_;
wire _2168_;
wire _2169_;
wire _2170_;
wire _2171_;
wire _2172_;
wire _2173_;
wire _2174_;
wire _2175_;
wire _2176_;
wire _2177_;
wire _2178_;
wire _2179_;
wire _2180_;
wire _2181_;
wire _2182_;
wire _2183_;
wire _2184_;
wire _2185_;
wire _2186_;
wire _2187_;
wire _2188_;
wire _2189_;
wire _2190_;
wire _2191_;
wire _2192_;
wire _2193_;
wire _2194_;
wire _2195_;
wire _2196_;
wire _2197_;
wire _2198_;
wire _2199_;
wire _2200_;
wire _2201_;
wire _2202_;
wire _2203_;
wire _2204_;
wire _2205_;
wire _2206_;
wire _2207_;
wire _2208_;
wire _2209_;
wire _2210_;
wire _2211_;
wire _2212_;
wire _2213_;
wire _2214_;
wire _2215_;
wire _2216_;
wire _2217_;
wire _2218_;
wire _2219_;
wire _2220_;
wire _2221_;
wire _2222_;
wire _2223_;
wire _2224_;
wire _2225_;
wire _2226_;
wire _2227_;
wire _2228_;
wire _2229_;
wire _2230_;
wire _2231_;
wire _2232_;
wire _2233_;
wire _2234_;
wire _2235_;
wire _2236_;
wire _2237_;
wire _2238_;
wire _2239_;
wire _2240_;
wire _2241_;
wire _2242_;
wire _2243_;
wire _2244_;
wire _2245_;
wire _2246_;
wire _2247_;
wire _2248_;
wire _2249_;
wire _2250_;
wire _2251_;
wire _2252_;
wire _2253_;
wire _2254_;
wire _2255_;
wire _2256_;
wire _2257_;
wire _2258_;
wire _2259_;
wire _2260_;
wire _2261_;
wire _2262_;
wire _2263_;
wire _2264_;
wire _2265_;
wire _2266_;
wire _2267_;
wire _2268_;
wire _2269_;
wire _2270_;
wire _2271_;
wire _2272_;
wire _2273_;
wire _2274_;
wire _2275_;
wire _2276_;
wire _2277_;
wire _2278_;
wire _2279_;
wire _2280_;
wire _2281_;
wire _2282_;
wire _2283_;
wire _2284_;
wire _2285_;
wire _2286_;
wire _2287_;
wire _2288_;
wire _2289_;
wire _2290_;
wire _2291_;
wire _2292_;
wire _2293_;
wire _2294_;
wire _2295_;
wire _2296_;
wire _2297_;
wire _2298_;
wire _2299_;
wire _2300_;
wire _2301_;
wire _2302_;
wire _2303_;
wire _2304_;
wire _2305_;
wire _2306_;
wire _2307_;
wire _2308_;
wire _2309_;
wire _2310_;
wire _2311_;
wire _2312_;
wire _2313_;
wire _2314_;
wire _2315_;
wire _2316_;
wire _2317_;
wire _2318_;
wire _2319_;
wire _2320_;
wire _2321_;
wire _2322_;
wire _2323_;
wire _2324_;
wire _2325_;
wire _2326_;
wire _2327_;
wire _2328_;
wire _2329_;
wire _2330_;
wire _2331_;
wire _2332_;
wire _2333_;
wire _2334_;
wire _2335_;
wire _2336_;
wire _2337_;
wire _2338_;
wire _2339_;
wire _2340_;
wire _2341_;
wire _2342_;
wire _2343_;
wire _2344_;
wire _2345_;
wire _2346_;
wire _2347_;
wire _2348_;
wire _2349_;
wire _2350_;
wire _2351_;
wire _2352_;
wire _2353_;
wire _2354_;
wire _2355_;
wire _2356_;
wire _2357_;
wire _2358_;
wire _2359_;
wire _2360_;
wire _2361_;
wire _2362_;
wire _2363_;
wire _2364_;
wire _2365_;
wire _2366_;
wire _2367_;
wire _2368_;
wire _2369_;
wire _2370_;
wire _2371_;
wire _2372_;
wire _2373_;
wire _2374_;
wire _2375_;
wire _2376_;
wire _2377_;
wire _2378_;
wire _2379_;
wire _2380_;
wire _2381_;
wire _2382_;
wire _2383_;
wire _2384_;
wire _2385_;
wire _2386_;
wire _2387_;
wire _2388_;
wire _2389_;
wire _2390_;
wire _2391_;
wire _2392_;
wire _2393_;
wire _2394_;
wire _2395_;
wire _2396_;
wire _2397_;
wire _2398_;
wire _2399_;
wire _2400_;
wire _2401_;
wire _2402_;
wire _2403_;
wire _2404_;
wire _2405_;
wire _2406_;
wire _2407_;
wire _2408_;
wire _2409_;
wire _2410_;
wire _2411_;
wire _2412_;
wire _2413_;
wire _2414_;
wire _2415_;
wire _2416_;
wire _2417_;
wire _2418_;
wire _2419_;
wire _2420_;
wire _2421_;
wire _2422_;
wire _2423_;
wire _2424_;
wire _2425_;
wire _2426_;
wire _2427_;
wire _2428_;
wire _2429_;
wire _2430_;
wire _2431_;
wire _2432_;
wire _2433_;
wire _2434_;
wire _2435_;
wire _2436_;
wire _2437_;
wire _2438_;
wire _2439_;
wire _2440_;
wire _2441_;
wire _2442_;
wire _2443_;
wire _2444_;
wire _2445_;
wire _2446_;
wire _2447_;
wire _2448_;
wire _2449_;
wire _2450_;
wire _2451_;
wire _2452_;
wire _2453_;
wire _2454_;
wire _2455_;
wire _2456_;
wire _2457_;
wire _2458_;
wire _2459_;
wire _2460_;
wire _2461_;
wire _2462_;
wire _2463_;
wire _2464_;
wire _2465_;
wire _2466_;
wire _2467_;
wire _2468_;
wire _2469_;
wire _2470_;
wire _2471_;
wire _2472_;
wire _2473_;
wire _2474_;
wire _2475_;
wire _2476_;
wire _2477_;
wire _2478_;
wire _2479_;
wire _2480_;
wire _2481_;
wire _2482_;
wire _2483_;
wire _2484_;
wire _2485_;
wire _2486_;
wire _2487_;
wire _2488_;
wire _2489_;
wire _2490_;
wire _2491_;
wire _2492_;
wire _2493_;
wire _2494_;
wire _2495_;
wire _2496_;
wire _2497_;
wire _2498_;
wire _2499_;
wire _2500_;
wire _2501_;
wire _2502_;
wire _2503_;
wire _2504_;
wire _2505_;
wire _2506_;
wire _2507_;
wire _2508_;
wire _2509_;
wire _2510_;
wire _2511_;
wire _2512_;
wire _2513_;
wire _2514_;
wire _2515_;
wire _2516_;
wire _2517_;
wire _2518_;
wire _2519_;
wire _2520_;
wire _2521_;
wire _2522_;
wire _2523_;
wire _2524_;
wire _2525_;
wire _2526_;
wire _2527_;
wire _2528_;
wire _2529_;
wire _2530_;
wire _2531_;
wire _2532_;
wire _2533_;
wire _2534_;
wire _2535_;
wire _2536_;
wire _2537_;
wire _2538_;
wire _2539_;
wire _2540_;
wire _2541_;
wire _2542_;
wire _2543_;
wire _2544_;
wire _2545_;
wire _2546_;
wire _2547_;
wire _2548_;
wire _2549_;
wire _2550_;
wire _2551_;
wire _2552_;
wire _2553_;
wire _2554_;
wire _2555_;
wire _2556_;
wire _2557_;
wire _2558_;
wire _2559_;
wire _2560_;
wire _2561_;
wire _2562_;
wire _2563_;
wire _2564_;
wire _2565_;
wire _2566_;
wire _2567_;
wire _2568_;
wire _2569_;
wire _2570_;
wire _2571_;
wire _2572_;
wire _2573_;
wire _2574_;
wire _2575_;
wire _2576_;
wire _2577_;
wire _2578_;
wire _2579_;
wire _2580_;
wire _2581_;
wire _2582_;
wire _2583_;
wire _2584_;
wire _2585_;
wire _2586_;
wire _2587_;
wire _2588_;
wire _2589_;
wire _2590_;
wire _2591_;
wire _2592_;
wire _2593_;
wire _2594_;
wire _2595_;
wire _2596_;
wire _2597_;
wire _2598_;
wire _2599_;
wire _2600_;
wire _2601_;
wire _2602_;
wire _2603_;
wire _2604_;
wire _2605_;
wire _2606_;
wire _2607_;
wire _2608_;
wire _2609_;
wire _2610_;
wire _2611_;
wire _2612_;
wire _2613_;
wire _2614_;
wire _2615_;
wire _2616_;
wire _2617_;
wire _2618_;
wire _2619_;
wire _2620_;
wire _2621_;
wire _2622_;
wire _2623_;
wire _2624_;
wire _2625_;
wire _2626_;
wire _2627_;
wire _2628_;
wire _2629_;
wire _2630_;
wire _2631_;
wire _2632_;
wire _2633_;
wire _2634_;
wire _2635_;
wire _2636_;
wire _2637_;
wire _2638_;
wire _2639_;
wire _2640_;
wire _2641_;
wire _2642_;
wire _2643_;
wire _2644_;
wire _2645_;
wire _2646_;
wire _2647_;
wire _2648_;
wire _2649_;
wire _2650_;
wire _2651_;
wire _2652_;
wire _2653_;
wire _2654_;
wire _2655_;
wire _2656_;
wire _2657_;
wire _2658_;
wire _2659_;
wire _2660_;
wire _2661_;
wire _2662_;
wire _2663_;
wire _2664_;
wire _2665_;
wire _2666_;
wire _2667_;
wire _2668_;
wire _2669_;
wire _2670_;
wire _2671_;
wire _2672_;
wire _2673_;
wire _2674_;
wire _2675_;
wire _2676_;
wire _2677_;
wire _2678_;
wire _2679_;
wire _2680_;
wire _2681_;
wire _2682_;
wire _2683_;
wire _2684_;
wire _2685_;
wire _2686_;
wire _2687_;
wire _2688_;
wire _2689_;
wire _2690_;
wire _2691_;
wire _2692_;
wire _2693_;
wire _2694_;
wire _2695_;
wire _2696_;
wire _2697_;
wire _2698_;
wire _2699_;
wire _2700_;
wire _2701_;
wire _2702_;
wire _2703_;
wire _2704_;
wire _2705_;
wire _2706_;
wire _2707_;
wire _2708_;
wire _2709_;
wire _2710_;
wire _2711_;
wire _2712_;
wire _2713_;
wire _2714_;
wire _2715_;
wire _2716_;
wire _2717_;
wire _2718_;
wire _2719_;
wire _2720_;
wire _2721_;
wire _2722_;
wire _2723_;
wire _2724_;
wire _2725_;
wire _2726_;
wire _2727_;
wire _2728_;
wire _2729_;
wire _2730_;
wire _2731_;
wire _2732_;
wire _2733_;
wire _2734_;
wire _2735_;
wire _2736_;
wire _2737_;
wire _2738_;
wire _2739_;
wire _2740_;
wire _2741_;
wire _2742_;
wire _2743_;
wire _2744_;
wire _2745_;
wire _2746_;
wire _2747_;
wire _2748_;
wire _2749_;
wire _2750_;
wire _2751_;
wire _2752_;
wire _2753_;
wire _2754_;
wire _2755_;
wire _2756_;
wire _2757_;
wire _2758_;
wire _2759_;
wire _2760_;
wire _2761_;
wire _2762_;
wire _2763_;
wire _2764_;
wire _2765_;
wire _2766_;
wire _2767_;
wire _2768_;
wire _2769_;
wire _2770_;
wire _2771_;
wire _2772_;
wire _2773_;
wire _2774_;
wire _2775_;
wire _2776_;
wire _2777_;
wire _2778_;
wire _2779_;
wire _2780_;
wire _2781_;
wire _2782_;
wire _2783_;
wire _2784_;
wire _2785_;
wire _2786_;
wire _2787_;
wire _2788_;
wire _2789_;
wire _2790_;
wire _2791_;
wire _2792_;
wire _2793_;
wire _2794_;
wire _2795_;
wire _2796_;
wire _2797_;
wire _2798_;
wire _2799_;
wire _2800_;
wire _2801_;
wire _2802_;
wire _2803_;
wire _2804_;
wire _2805_;
wire _2806_;
wire _2807_;
wire _2808_;
wire _2809_;
wire _2810_;
wire _2811_;
wire _2812_;
wire _2813_;
wire _2814_;
wire _2815_;
wire _2816_;
wire _2817_;
wire _2818_;
wire _2819_;
wire _2820_;
wire _2821_;
wire _2822_;
wire _2823_;
wire _2824_;
wire _2825_;
wire _2826_;
wire _2827_;
wire _2828_;
wire _2829_;
wire _2830_;
wire _2831_;
wire _2832_;
wire _2833_;
wire _2834_;
wire _2835_;
wire _2836_;
wire _2837_;
wire _2838_;
wire _2839_;
wire _2840_;
wire _2841_;
wire _2842_;
wire _2843_;
wire _2844_;
wire _2845_;
wire _2846_;
wire _2847_;
wire _2848_;
wire _2849_;
wire _2850_;
wire _2851_;
wire _2852_;
wire _2853_;
wire _2854_;
wire _2855_;
wire _2856_;
wire _2857_;
wire _2858_;
wire _2859_;
wire _2860_;
wire _2861_;
wire _2862_;
wire _2863_;
wire _2864_;
wire _2865_;
wire _2866_;
wire _2867_;
wire _2868_;
wire _2869_;
wire _2870_;
wire _2871_;
wire _2872_;
wire _2873_;
wire _2874_;
wire _2875_;
wire _2876_;
wire _2877_;
wire _2878_;
wire _2879_;
wire _2880_;
wire _2881_;
wire _2882_;
wire _2883_;
wire _2884_;
wire _2885_;
wire _2886_;
wire _2887_;
wire _2888_;
wire _2889_;
wire _2890_;
wire _2891_;
wire _2892_;
wire _2893_;
wire _2894_;
wire _2895_;
wire _2896_;
wire _2897_;
wire _2898_;
wire _2899_;
wire _2900_;
wire _2901_;
wire _2902_;
wire _2903_;
wire _2904_;
wire _2905_;
wire _2906_;
wire _2907_;
wire _2908_;
wire _2909_;
wire _2910_;
wire _2911_;
wire _2912_;
wire _2913_;
wire _2914_;
wire _2915_;
wire _2916_;
wire _2917_;
wire _2918_;
wire _2919_;
wire _2920_;
wire _2921_;
wire _2922_;
wire _2923_;
wire _2924_;
wire _2925_;
wire _2926_;
wire _2927_;
wire _2928_;
wire _2929_;
wire _2930_;
wire _2931_;
wire _2932_;
wire _2933_;
wire _2934_;
wire _2935_;
wire _2936_;
wire _2937_;
wire _2938_;
wire _2939_;
wire _2940_;
wire _2941_;
wire _2942_;
wire _2943_;
wire _2944_;
wire _2945_;
wire _2946_;
wire _2947_;
wire _2948_;
wire _2949_;
wire _2950_;
wire _2951_;
wire _2952_;
wire _2953_;
wire _2954_;
wire _2955_;
wire _2956_;
wire _2957_;
wire _2958_;
wire _2959_;
wire _2960_;
wire _2961_;
wire _2962_;
wire _2963_;
wire _2964_;
wire _2965_;
wire _2966_;
wire _2967_;
wire _2968_;
wire _2969_;
wire _2970_;
wire _2971_;
wire _2972_;
wire _2973_;
wire _2974_;
wire _2975_;
wire _2976_;
wire _2977_;
wire _2978_;
wire _2979_;
wire _2980_;
wire _2981_;
wire _2982_;
wire _2983_;
wire _2984_;
wire _2985_;
wire _2986_;
wire _2987_;
wire _2988_;
wire _2989_;
wire _2990_;
wire _2991_;
wire _2992_;
wire _2993_;
wire _2994_;
wire _2995_;
wire _2996_;
wire _2997_;
wire _2998_;
wire _2999_;
wire _3000_;
wire _3001_;
wire _3002_;
wire _3003_;
wire _3004_;
wire _3005_;
wire _3006_;
wire _3007_;
wire _3008_;
wire _3009_;
wire _3010_;
wire _3011_;
wire _3012_;
wire _3013_;
wire _3014_;
wire _3015_;
wire _3016_;
wire _3017_;
wire _3018_;
wire _3019_;
wire _3020_;
wire _3021_;
wire _3022_;
wire _3023_;
wire _3024_;
wire _3025_;
wire _3026_;
wire _3027_;
wire _3028_;
wire _3029_;
wire _3030_;
wire _3031_;
wire _3032_;
wire _3033_;
wire _3034_;
wire _3035_;
wire _3036_;
wire _3037_;
wire _3038_;
wire _3039_;
wire _3040_;
wire _3041_;
wire _3042_;
wire _3043_;
wire _3044_;
wire _3045_;
wire _3046_;
wire _3047_;
wire _3048_;
wire _3049_;
wire _3050_;
wire _3051_;
wire _3052_;
wire _3053_;
wire _3054_;
wire _3055_;
wire _3056_;
wire _3057_;
wire _3058_;
wire _3059_;
wire _3060_;
wire _3061_;
wire _3062_;
wire _3063_;
wire _3064_;
wire _3065_;
wire _3066_;
wire _3067_;
wire _3068_;
wire _3069_;
wire _3070_;
wire _3071_;
wire _3072_;
wire _3073_;
wire _3074_;
wire _3075_;
wire _3076_;
wire _3077_;
wire _3078_;
wire _3079_;
wire _3080_;
wire _3081_;
wire _3082_;
wire _3083_;
wire _3084_;
wire _3085_;
wire _3086_;
wire _3087_;
wire _3088_;
wire _3089_;
wire _3090_;
wire _3091_;
wire _3092_;
wire _3093_;
wire _3094_;
wire _3095_;
wire _3096_;
wire _3097_;
wire _3098_;
wire _3099_;
wire _3100_;
wire _3101_;
wire _3102_;
wire _3103_;
wire _3104_;
wire _3105_;
wire _3106_;
wire _3107_;
wire _3108_;
wire _3109_;
wire _3110_;
wire _3111_;
wire _3112_;
wire _3113_;
wire _3114_;
wire _3115_;
wire _3116_;
wire _3117_;
wire _3118_;
wire _3119_;
wire _3120_;
wire _3121_;
wire _3122_;
wire _3123_;
wire _3124_;
wire _3125_;
wire _3126_;
wire _3127_;
wire _3128_;
wire _3129_;
wire _3130_;
wire _3131_;
wire _3132_;
wire _3133_;
wire _3134_;
wire _3135_;
wire _3136_;
wire _3137_;
wire _3138_;
wire _3139_;
wire _3140_;
wire _3141_;
wire _3142_;
wire _3143_;
wire _3144_;
wire _3145_;
wire _3146_;
wire _3147_;
wire _3148_;
wire _3149_;
wire _3150_;
wire _3151_;
wire _3152_;
wire _3153_;
wire _3154_;
wire _3155_;
wire _3156_;
wire _3157_;
wire _3158_;
wire _3159_;
wire _3160_;
wire _3161_;
wire _3162_;
wire _3163_;
wire _3164_;
wire _3165_;
wire _3166_;
wire _3167_;
wire _3168_;
wire _3169_;
wire _3170_;
wire _3171_;
wire _3172_;
wire _3173_;
wire _3174_;
wire _3175_;
wire _3176_;
wire _3177_;
wire _3178_;
wire _3179_;
wire _3180_;
wire _3181_;
wire _3182_;
wire _3183_;
wire _3184_;
wire _3185_;
wire _3186_;
wire _3187_;
wire _3188_;
wire _3189_;
wire _3190_;
wire _3191_;
wire _3192_;
wire _3193_;
wire _3194_;
wire _3195_;
wire _3196_;
wire _3197_;
wire _3198_;
wire _3199_;
wire _3200_;
wire _3201_;
wire _3202_;
wire _3203_;
wire _3204_;
wire _3205_;
wire _3206_;
wire _3207_;
wire _3208_;
wire _3209_;
wire _3210_;
wire _3211_;
wire _3212_;
wire _3213_;
wire _3214_;
wire _3215_;
wire _3216_;
wire _3217_;
wire _3218_;
wire _3219_;
wire _3220_;
wire _3221_;
wire _3222_;
wire _3223_;
wire _3224_;
wire _3225_;
wire _3226_;
wire _3227_;
wire _3228_;
wire _3229_;
wire _3230_;
wire _3231_;
wire _3232_;
wire _3233_;
wire _3234_;
wire _3235_;
wire _3236_;
wire _3237_;
wire _3238_;
wire _3239_;
wire _3240_;
wire _3241_;
wire _3242_;
wire _3243_;
wire _3244_;
wire _3245_;
wire _3246_;
wire _3247_;
wire _3248_;
wire _3249_;
wire _3250_;
wire _3251_;
wire _3252_;
wire _3253_;
wire _3254_;
wire _3255_;
wire _3256_;
wire _3257_;
wire _3258_;
wire _3259_;
wire _3260_;
wire _3261_;
wire _3262_;
wire _3263_;
wire _3264_;
wire _3265_;
wire _3266_;
wire _3267_;
wire _3268_;
wire _3269_;
wire _3270_;
wire _3271_;
wire _3272_;
wire _3273_;
wire _3274_;
wire _3275_;
wire _3276_;
wire _3277_;
wire _3278_;
wire _3279_;
wire _3280_;
wire _3281_;
wire _3282_;
wire _3283_;
wire _3284_;
wire _3285_;
wire _3286_;
wire _3287_;
wire _3288_;
wire _3289_;
wire _3290_;
wire _3291_;
wire _3292_;
wire _3293_;
wire _3294_;
wire _3295_;
wire _3296_;
wire _3297_;
wire _3298_;
wire _3299_;
wire _3300_;
wire _3301_;
wire _3302_;
wire _3303_;
wire _3304_;
wire _3305_;
wire _3306_;
wire _3307_;
wire _3308_;
wire _3309_;
wire _3310_;
wire _3311_;
wire _3312_;
wire _3313_;
wire _3314_;
wire _3315_;
wire _3316_;
wire _3317_;
wire _3318_;
wire _3319_;
wire _3320_;
wire _3321_;
wire _3322_;
wire _3323_;
wire _3324_;
wire _3325_;
wire _3326_;
wire _3327_;
wire _3328_;
wire _3329_;
wire _3330_;
wire _3331_;
wire _3332_;
wire _3333_;
wire _3334_;
wire _3335_;
wire _3336_;
wire _3337_;
wire _3338_;
wire _3339_;
wire _3340_;
wire _3341_;
wire _3342_;
wire _3343_;
wire _3344_;
wire _3345_;
wire _3346_;
wire _3347_;
wire _3348_;
wire _3349_;
wire _3350_;
wire _3351_;
wire _3352_;
wire _3353_;
wire _3354_;
wire _3355_;
wire _3356_;
wire _3357_;
wire _3358_;
wire _3359_;
wire _3360_;
wire _3361_;
wire _3362_;
wire _3363_;
wire _3364_;
wire _3365_;
wire _3366_;
wire _3367_;
wire _3368_;
wire _3369_;
wire _3370_;
wire _3371_;
wire _3372_;
wire _3373_;
wire _3374_;
wire _3375_;
wire _3376_;
wire _3377_;
wire _3378_;
wire _3379_;
wire _3380_;
wire _3381_;
wire _3382_;
wire _3383_;
wire _3384_;
wire _3385_;
wire _3386_;
wire _3387_;
wire _3388_;
wire _3389_;
wire _3390_;
wire _3391_;
wire _3392_;
wire _3393_;
wire _3394_;
wire _3395_;
wire _3396_;
wire _3397_;
wire _3398_;
wire _3399_;
wire _3400_;
wire _3401_;
wire _3402_;
wire _3403_;
wire _3404_;
wire _3405_;
wire _3406_;
wire _3407_;
wire _3408_;
wire _3409_;
wire _3410_;
wire _3411_;
wire _3412_;
wire _3413_;
wire _3414_;
wire _3415_;
wire _3416_;
wire _3417_;
wire _3418_;
wire _3419_;
wire _3420_;
wire _3421_;
wire _3422_;
wire _3423_;
wire _3424_;
wire _3425_;
wire _3426_;
wire _3427_;
wire _3428_;
wire _3429_;
wire _3430_;
wire _3431_;
wire _3432_;
wire _3433_;
wire _3434_;
wire _3435_;
wire _3436_;
wire _3437_;
wire _3438_;
wire _3439_;
wire _3440_;
wire _3441_;
wire _3442_;
wire _3443_;
wire _3444_;
wire _3445_;
wire _3446_;
wire _3447_;
wire _3448_;
wire _3449_;
wire _3450_;
wire _3451_;
wire _3452_;
wire _3453_;
wire _3454_;
wire _3455_;
wire _3456_;
wire _3457_;
wire _3458_;
wire _3459_;
wire _3460_;
wire _3461_;
wire _3462_;
wire _3463_;
wire _3464_;
wire _3465_;
wire _3466_;
wire _3467_;
wire _3468_;
wire _3469_;
wire _3470_;
wire _3471_;
wire _3472_;
wire _3473_;
wire _3474_;
wire _3475_;
wire _3476_;
wire _3477_;
wire _3478_;
wire _3479_;
wire _3480_;
wire _3481_;
wire _3482_;
wire _3483_;
wire _3484_;
wire _3485_;
wire _3486_;
wire _3487_;
wire _3488_;
wire _3489_;
wire _3490_;
wire _3491_;
wire _3492_;
wire _3493_;
wire _3494_;
wire _3495_;
wire _3496_;
wire _3497_;
wire _3498_;
wire _3499_;
wire _3500_;
wire _3501_;
wire _3502_;
wire _3503_;
wire _3504_;
wire _3505_;
wire _3506_;
wire _3507_;
wire _3508_;
wire _3509_;
wire _3510_;
wire _3511_;
wire _3512_;
wire _3513_;
wire _3514_;
wire _3515_;
wire _3516_;
wire _3517_;
wire _3518_;
wire _3519_;
wire _3520_;
wire _3521_;
wire _3522_;
wire _3523_;
wire _3524_;
wire _3525_;
wire _3526_;
wire _3527_;
wire _3528_;
wire _3529_;
wire _3530_;
wire _3531_;
wire _3532_;
wire _3533_;
wire _3534_;
wire _3535_;
wire _3536_;
wire _3537_;
wire _3538_;
wire _3539_;
wire _3540_;
wire _3541_;
wire _3542_;
wire _3543_;
wire _3544_;
wire _3545_;
wire _3546_;
wire _3547_;
wire _3548_;
wire _3549_;
wire _3550_;
wire _3551_;
wire _3552_;
wire _3553_;
wire _3554_;
wire _3555_;
wire _3556_;
wire _3557_;
wire _3558_;
wire _3559_;
wire _3560_;
wire _3561_;
wire _3562_;
wire _3563_;
wire _3564_;
wire _3565_;
wire _3566_;
wire _3567_;
wire _3568_;
wire _3569_;
wire _3570_;
wire _3571_;
wire _3572_;
wire _3573_;
wire _3574_;
wire _3575_;
wire _3576_;
wire _3577_;
wire _3578_;
wire _3579_;
wire _3580_;
wire _3581_;
wire _3582_;
wire _3583_;
wire _3584_;
wire _3585_;
wire _3586_;
wire _3587_;
wire _3588_;
wire _3589_;
wire _3590_;
wire _3591_;
wire _3592_;
wire _3593_;
wire _3594_;
wire _3595_;
wire _3596_;
wire _3597_;
wire _3598_;
wire _3599_;
wire _3600_;
wire _3601_;
wire _3602_;
wire _3603_;
wire _3604_;
wire _3605_;
wire _3606_;
wire _3607_;
wire _3608_;
wire _3609_;
wire _3610_;
wire _3611_;
wire _3612_;
wire _3613_;
wire _3614_;
wire _3615_;
wire _3616_;
wire _3617_;
wire _3618_;
wire _3619_;
wire _3620_;
wire _3621_;
wire _3622_;
wire _3623_;
wire _3624_;
wire _3625_;
wire _3626_;
wire _3627_;
wire _3628_;
wire _3629_;
wire _3630_;
wire _3631_;
wire _3632_;
wire _3633_;
wire _3634_;
wire _3635_;
wire _3636_;
wire _3637_;
wire _3638_;
wire _3639_;
wire _3640_;
wire _3641_;
wire _3642_;
wire _3643_;
wire _3644_;
wire _3645_;
wire _3646_;
wire _3647_;
wire _3648_;
wire _3649_;
wire _3650_;
wire _3651_;
wire _3652_;
wire _3653_;
wire _3654_;
wire _3655_;
wire _3656_;
wire _3657_;
wire _3658_;
wire _3659_;
wire _3660_;
wire _3661_;
wire _3662_;
wire _3663_;
wire _3664_;
wire _3665_;
wire _3666_;
wire _3667_;
wire _3668_;
wire _3669_;
wire _3670_;
wire _3671_;
wire _3672_;
wire _3673_;
wire _3674_;
wire _3675_;
wire _3676_;
wire _3677_;
wire _3678_;
wire _3679_;
wire _3680_;
wire _3681_;
wire _3682_;
wire _3683_;
wire _3684_;
wire _3685_;
wire _3686_;
wire _3687_;
wire _3688_;
wire _3689_;
wire _3690_;
wire _3691_;
wire _3692_;
wire _3693_;
wire _3694_;
wire _3695_;
wire _3696_;
wire _3697_;
wire _3698_;
wire _3699_;
wire _3700_;
wire _3701_;
wire _3702_;
wire _3703_;
wire _3704_;
wire _3705_;
wire _3706_;
wire _3707_;
wire _3708_;
wire _3709_;
wire _3710_;
wire _3711_;
wire _3712_;
wire _3713_;
wire _3714_;
wire _3715_;
wire _3716_;
wire _3717_;
wire _3718_;
wire _3719_;
wire _3720_;
wire _3721_;
wire _3722_;
wire _3723_;
wire _3724_;
wire _3725_;
wire _3726_;
wire _3727_;
wire _3728_;
wire _3729_;
wire _3730_;
wire _3731_;
wire _3732_;
wire _3733_;
wire _3734_;
wire _3735_;
wire _3736_;
wire _3737_;
wire _3738_;
wire _3739_;
wire _3740_;
wire _3741_;
wire _3742_;
wire _3743_;
wire _3744_;
wire _3745_;
wire _3746_;
wire _3747_;
wire _3748_;
wire _3749_;
wire _3750_;
wire _3751_;
wire _3752_;
wire _3753_;
wire _3754_;
wire _3755_;
wire _3756_;
wire _3757_;
wire _3758_;
wire _3759_;
wire _3760_;
wire _3761_;
wire _3762_;
wire _3763_;
wire _3764_;
wire _3765_;
wire _3766_;
wire _3767_;
wire _3768_;
wire _3769_;
wire _3770_;
wire _3771_;
wire _3772_;
wire _3773_;
wire _3774_;
wire _3775_;
wire _3776_;
wire _3777_;
wire _3778_;
wire _3779_;
wire _3780_;
wire _3781_;
wire _3782_;
wire _3783_;
wire _3784_;
wire _3785_;
wire _3786_;
wire _3787_;
wire _3788_;
wire _3789_;
wire _3790_;
wire _3791_;
wire _3792_;
wire _3793_;
wire _3794_;
wire _3795_;
wire _3796_;
wire _3797_;
wire _3798_;
wire _3799_;
wire _3800_;
wire _3801_;
wire _3802_;
wire _3803_;
wire _3804_;
wire _3805_;
wire _3806_;
wire _3807_;
wire _3808_;
wire _3809_;
wire _3810_;
wire _3811_;
wire _3812_;
wire _3813_;
wire _3814_;
wire _3815_;
wire _3816_;
wire _3817_;
wire _3818_;
wire _3819_;
wire _3820_;
wire _3821_;
wire _3822_;
wire _3823_;
wire _3824_;
wire _3825_;
wire _3826_;
wire _3827_;
wire _3828_;
wire _3829_;
wire _3830_;
wire _3831_;
wire _3832_;
wire _3833_;
wire _3834_;
wire _3835_;
wire _3836_;
wire _3837_;
wire _3838_;
wire _3839_;
wire _3840_;
wire _3841_;
wire _3842_;
wire _3843_;
wire _3844_;
wire _3845_;
wire _3846_;
wire _3847_;
wire _3848_;
wire _3849_;
wire _3850_;
wire _3851_;
wire _3852_;
wire _3853_;
wire _3854_;
wire _3855_;
wire _3856_;
wire _3857_;
wire _3858_;
wire _3859_;
wire _3860_;
wire _3861_;
wire _3862_;
wire _3863_;
wire _3864_;
wire _3865_;
wire _3866_;
wire _3867_;
wire _3868_;
wire _3869_;
wire _3870_;
wire _3871_;
wire _3872_;
wire _3873_;
wire _3874_;
wire _3875_;
wire _3876_;
wire _3877_;
wire _3878_;
wire _3879_;
wire _3880_;
wire _3881_;
wire _3882_;
wire _3883_;
wire _3884_;
wire _3885_;
wire _3886_;
wire _3887_;
wire _3888_;
wire _3889_;
wire _3890_;
wire _3891_;
wire _3892_;
wire _3893_;
wire _3894_;
wire _3895_;
wire _3896_;
wire _3897_;
wire _3898_;
wire _3899_;
wire _3900_;
wire _3901_;
wire _3902_;
wire _3903_;
wire _3904_;
wire _3905_;
wire _3906_;
wire _3907_;
wire _3908_;
wire _3909_;
wire _3910_;
wire _3911_;
wire _3912_;
wire _3913_;
wire _3914_;
wire _3915_;
wire _3916_;
wire _3917_;
wire _3918_;
wire _3919_;
wire _3920_;
wire _3921_;
wire _3922_;
wire _3923_;
wire _3924_;
wire _3925_;
wire _3926_;
wire _3927_;
wire _3928_;
wire _3929_;
wire _3930_;
wire _3931_;
wire _3932_;
wire _3933_;
wire _3934_;
wire _3935_;
wire _3936_;
wire _3937_;
wire _3938_;
wire _3939_;
wire _3940_;
wire _3941_;
wire _3942_;
wire _3943_;
wire _3944_;
wire _3945_;
wire _3946_;
wire _3947_;
wire _3948_;
wire _3949_;
wire _3950_;
wire _3951_;
wire _3952_;
wire _3991_;
wire _3992_;
wire _3993_;
wire _3994_;
wire _3995_;
wire _3996_;
wire _3997_;
wire _3998_;
wire _3999_;
wire _4000_;
wire _4001_;
wire _4002_;
wire _4003_;
wire _4008_;
wire _4009_;
wire _4010_;
wire _4011_;
wire _4012_;
wire _4013_;
wire _4014_;
wire _4015_;
wire _4016_;
wire _4017_;
wire _4018_;
wire _4019_;
wire _4020_;
wire _4021_;
wire _4022_;
wire _4023_;
wire _4024_;
wire _4025_;
wire _4026_;
wire _4027_;
wire _4028_;
wire _4029_;
wire _4042_;
wire _4043_;
wire _4044_;
wire _4045_;
wire _4046_;
wire _4047_;
wire _4048_;
wire _4049_;
wire _4050_;
wire _4051_;
wire _4052_;
wire _4053_;
wire _4054_;
wire _4055_;
wire _4056_;
wire _4057_;
wire _4058_;
wire _4059_;
wire _4060_;
wire _4061_;
wire _4062_;
wire _4063_;
wire _4064_;
wire _4065_;
wire _4066_;
wire _4067_;
wire _4068_;
wire _4069_;
wire _4070_;
wire _4071_;
wire _4072_;
wire _4073_;
wire _4074_;
wire _4075_;
wire _4076_;
wire _4077_;
wire _4078_;
wire _4079_;
wire _4080_;
wire _4081_;
wire _4082_;
wire _4083_;
wire _4084_;
wire _4085_;
wire _4086_;
wire _4087_;
wire _4088_;
wire _4089_;
wire _4090_;
wire _4091_;
wire _4092_;
wire _4093_;
wire _4094_;
wire _4095_;
wire _4096_;
wire _4097_;
wire _4098_;
wire _4099_;
wire _4100_;
wire _4101_;
wire _4102_;
wire _4103_;
wire _4104_;
wire _4105_;
wire _4106_;
wire _4107_;
wire _4108_;
wire _4109_;
wire _4110_;
wire _4111_;
wire _4112_;
wire _4113_;
wire _4114_;
wire _4115_;
wire _4116_;
wire _4117_;
wire _4118_;
wire _4119_;
wire _4120_;
wire _4121_;
wire _4122_;
wire _4123_;
wire _4144_;
wire _4145_;
wire _4146_;
wire _4147_;
wire _4148_;
wire _4149_;
wire _4150_;
wire _4151_;
wire _4152_;
wire _4153_;
wire _4154_;
wire _4155_;
wire _4156_;
wire _4157_;
wire _4158_;
wire _4159_;
wire _4160_;
wire _4161_;
wire _4162_;
wire _4163_;
wire _4164_;
wire _4165_;
wire _4166_;
wire _4167_;
wire _4168_;
wire _4169_;
wire _4170_;
wire _4171_;
wire _4172_;
wire _4173_;
wire _4174_;
wire _4175_;
wire _4176_;
wire _4177_;
wire _4178_;
wire _4179_;
wire _4180_;
wire _4181_;
wire _4182_;
wire _4183_;
wire _4184_;
wire _4185_;
wire _4186_;
wire _4187_;
wire _4188_;
wire _4189_;
wire _4190_;
wire _4191_;
wire _4192_;
wire _4193_;
wire _4194_;
wire _4195_;
wire _4196_;
wire _4197_;
wire _4198_;
wire _4199_;
wire _4200_;
wire _4201_;
wire _4202_;
wire _4203_;
wire _4204_;
wire _4205_;
wire _4206_;
wire _4207_;
wire _4208_;
wire _4209_;
wire _4210_;
wire _4211_;
wire _4212_;
wire _4213_;
wire _4214_;
wire _4215_;
wire _4216_;
wire _4217_;
wire _4218_;
wire _4219_;
wire _4220_;
wire _4221_;
wire _4222_;
wire _4223_;
wire _4224_;
wire _4225_;
wire _4226_;
wire _4227_;
wire _4228_;
wire _4229_;
wire _4230_;
wire _4231_;
wire _4232_;
wire _4233_;
wire _4234_;
wire _4235_;
wire _4236_;
wire _4237_;
wire _4238_;
wire _4239_;
wire _4240_;
wire _4241_;
wire _4242_;
wire _4243_;
wire _4244_;
wire _4245_;
wire _4246_;
wire _4247_;
wire _4248_;
wire _4249_;
wire _4250_;
wire _4251_;
wire _4252_;
wire _4253_;
wire _4254_;
wire _4255_;
wire _4256_;
wire _4257_;
wire _4258_;
wire _4259_;
wire _4260_;
wire _4261_;
wire _4262_;
wire _4263_;
wire _4264_;
wire _4265_;
wire _4266_;
wire _4267_;
wire _4268_;
wire _4269_;
wire _4270_;
wire _4271_;
wire _4272_;
wire _4273_;
wire _4274_;
wire _4275_;
wire _4276_;
wire _4277_;
wire _4278_;
wire _4279_;
wire _4280_;
wire _4281_;
wire _4282_;
wire _4283_;
wire _4284_;
wire _4285_;
wire _4286_;
wire _4287_;
wire _4288_;
wire _4291_;
wire _4292_;
wire _4293_;
wire _4294_;
wire _4295_;
wire _4296_;
wire _4297_;
wire _4298_;
wire _4299_;
wire _4300_;
wire _4301_;
wire _4302_;
wire _4303_;
wire _4304_;
wire _4305_;
wire _4306_;
wire _4307_;
wire _4308_;
wire _4309_;
wire _4310_;
wire _4311_;
wire _4312_;
wire _4313_;
wire _4314_;
wire _4315_;
wire _4316_;
wire _4317_;
wire _4318_;
wire _4319_;
wire _4320_;
wire _4321_;
wire _4322_;
wire _4323_;
wire _4324_;
wire _4325_;
wire _4326_;
wire _4327_;
wire _4328_;
wire _4329_;
wire _4330_;
wire _4331_;
wire _4332_;
wire _4333_;
wire _4334_;
wire _4335_;
wire _4336_;
wire _4337_;
wire _4338_;
wire _4339_;
wire _4340_;
wire _4341_;
wire _4342_;
wire _4343_;
wire _4344_;
wire _4345_;
wire _4346_;
wire _4347_;
wire _4348_;
wire _4349_;
wire _4350_;
wire _4351_;
wire _4352_;
wire _4353_;
wire _4354_;
wire _4355_;
wire _4356_;
wire _4357_;
wire _4358_;
wire _4359_;
wire _4360_;
wire _4361_;
wire _4362_;
wire _4363_;
wire _4364_;
wire _4365_;
wire _4366_;
wire _4367_;
wire _4368_;
wire _4369_;
wire _4370_;
wire _4371_;
wire _4372_;
wire _4373_;
wire _4374_;
wire _4375_;
wire _4376_;
wire _4377_;
wire _4378_;
wire _4379_;
wire _4380_;
wire _4381_;
wire _4382_;
wire _4383_;
wire _4384_;
wire _4385_;
wire _4386_;
wire _4387_;
wire _4388_;
wire _4389_;
wire _4390_;
wire _4391_;
wire _4392_;
wire _4393_;
wire _4394_;
wire _4395_;
wire _4396_;
wire _4397_;
wire _4398_;
wire _4399_;
wire _4400_;
wire _4401_;
wire _4402_;
wire _4403_;
wire _4404_;
wire _4405_;
wire _4406_;
wire _4407_;
wire _4408_;
wire _4409_;
wire _4410_;
wire _4411_;
wire _4412_;
wire _4413_;
wire _4414_;
wire _4415_;
wire _4416_;
wire _4417_;
wire _4418_;
wire _4419_;
wire _4420_;
wire _4421_;
wire _4422_;
wire _4423_;
wire _4424_;
wire _4425_;
wire _4426_;
wire _4427_;
wire _4428_;
wire _4429_;
wire _4430_;
wire _4431_;
wire _4432_;
wire _4433_;
wire _4434_;
wire _4435_;
wire _4436_;
wire _4437_;
wire _4438_;
wire _4439_;
wire _4440_;
wire _4441_;
wire _4442_;
wire _4443_;
wire _4444_;
wire _4445_;
wire _4446_;
wire _4447_;
wire _4448_;
wire _4449_;
wire _4450_;
wire _4451_;
wire _4452_;
wire _4453_;
wire _4454_;
wire _4455_;
wire _4456_;
wire _4457_;
wire _4458_;
wire _4459_;
wire _4460_;
wire _4461_;
wire _4462_;
wire _4463_;
wire _4464_;
wire _4465_;
wire _4466_;
wire _4467_;
wire _4468_;
wire _4469_;
wire _4470_;
wire _4471_;
wire _4472_;
wire _4473_;
wire _4474_;
wire _4475_;
wire _4476_;
wire _4477_;
wire _4478_;
wire _4479_;
wire _4480_;
wire _4481_;
wire _4482_;
wire _4483_;
wire _4484_;
wire _4485_;
wire _4486_;
wire _4487_;
wire _4488_;
wire _4489_;
wire _4490_;
wire _4491_;
wire _4492_;
wire _4493_;
wire _4494_;
wire _4495_;
wire _4496_;
wire _4497_;
wire _4498_;
wire _4499_;
wire _4500_;
wire _4501_;
wire _4502_;
wire _4503_;
wire _4504_;
wire _4505_;
wire _4506_;
wire _4507_;
wire _4508_;
wire _4509_;
wire _4510_;
wire _4511_;
wire _4512_;
wire _4513_;
wire _4514_;
wire _4515_;
wire _4516_;
wire _4517_;
wire _4518_;
wire _4519_;
wire _4520_;
wire _4521_;
wire _4522_;
wire _4523_;
wire _4524_;
wire _4525_;
wire _4526_;
wire _4527_;
wire _4528_;
wire _4529_;
wire _4530_;
wire _4531_;
wire _4532_;
wire _4533_;
wire _4534_;
wire _4535_;
wire _4536_;
wire _4537_;
wire _4538_;
wire _4539_;
wire _4540_;
wire _4541_;
wire _4542_;
wire _4543_;
wire _4544_;
wire _4545_;
wire _4546_;
wire _4547_;
wire _4548_;
wire _4549_;
wire _4550_;
wire _4551_;
wire _4552_;
wire _4553_;
wire _4554_;
wire _4555_;
wire _4556_;
wire _4557_;
wire _4558_;
wire _4559_;
wire _4560_;
wire _4561_;
wire _4562_;
wire _4563_;
wire _4564_;
wire _4565_;
wire _4566_;
wire _4567_;
wire _4568_;
wire _4569_;
wire _4570_;
wire _4571_;
wire _4572_;
wire \d_pipe[10][12] ;
wire \d_pipe[10][13] ;
wire \d_pipe[10][14] ;
wire \d_pipe[10][15] ;
wire \d_pipe[10][16] ;
wire \d_pipe[10][17] ;
wire \d_pipe[10][18] ;
wire \d_pipe[10][19] ;
wire \d_pipe[10][20] ;
wire \d_pipe[10][21] ;
wire \d_pipe[10][22] ;
wire \d_pipe[10][23] ;
wire \d_pipe[11][12] ;
wire \d_pipe[11][13] ;
wire \d_pipe[11][14] ;
wire \d_pipe[11][15] ;
wire \d_pipe[11][16] ;
wire \d_pipe[11][17] ;
wire \d_pipe[11][18] ;
wire \d_pipe[11][19] ;
wire \d_pipe[11][20] ;
wire \d_pipe[11][21] ;
wire \d_pipe[11][22] ;
wire \d_pipe[11][23] ;
wire \d_pipe[1][12] ;
wire \d_pipe[1][13] ;
wire \d_pipe[1][14] ;
wire \d_pipe[1][15] ;
wire \d_pipe[1][16] ;
wire \d_pipe[1][17] ;
wire \d_pipe[1][18] ;
wire \d_pipe[1][19] ;
wire \d_pipe[1][20] ;
wire \d_pipe[1][21] ;
wire \d_pipe[1][22] ;
wire \d_pipe[1][23] ;
wire \d_pipe[2][12] ;
wire \d_pipe[2][13] ;
wire \d_pipe[2][14] ;
wire \d_pipe[2][15] ;
wire \d_pipe[2][16] ;
wire \d_pipe[2][17] ;
wire \d_pipe[2][18] ;
wire \d_pipe[2][19] ;
wire \d_pipe[2][20] ;
wire \d_pipe[2][21] ;
wire \d_pipe[2][22] ;
wire \d_pipe[2][23] ;
wire \d_pipe[3][12] ;
wire \d_pipe[3][13] ;
wire \d_pipe[3][14] ;
wire \d_pipe[3][15] ;
wire \d_pipe[3][16] ;
wire \d_pipe[3][17] ;
wire \d_pipe[3][18] ;
wire \d_pipe[3][19] ;
wire \d_pipe[3][20] ;
wire \d_pipe[3][21] ;
wire \d_pipe[3][22] ;
wire \d_pipe[3][23] ;
wire \d_pipe[4][12] ;
wire \d_pipe[4][13] ;
wire \d_pipe[4][14] ;
wire \d_pipe[4][15] ;
wire \d_pipe[4][16] ;
wire \d_pipe[4][17] ;
wire \d_pipe[4][18] ;
wire \d_pipe[4][19] ;
wire \d_pipe[4][20] ;
wire \d_pipe[4][21] ;
wire \d_pipe[4][22] ;
wire \d_pipe[4][23] ;
wire \d_pipe[5][12] ;
wire \d_pipe[5][13] ;
wire \d_pipe[5][14] ;
wire \d_pipe[5][15] ;
wire \d_pipe[5][16] ;
wire \d_pipe[5][17] ;
wire \d_pipe[5][18] ;
wire \d_pipe[5][19] ;
wire \d_pipe[5][20] ;
wire \d_pipe[5][21] ;
wire \d_pipe[5][22] ;
wire \d_pipe[5][23] ;
wire \d_pipe[6][12] ;
wire \d_pipe[6][13] ;
wire \d_pipe[6][14] ;
wire \d_pipe[6][15] ;
wire \d_pipe[6][16] ;
wire \d_pipe[6][17] ;
wire \d_pipe[6][18] ;
wire \d_pipe[6][19] ;
wire \d_pipe[6][20] ;
wire \d_pipe[6][21] ;
wire \d_pipe[6][22] ;
wire \d_pipe[6][23] ;
wire \d_pipe[7][12] ;
wire \d_pipe[7][13] ;
wire \d_pipe[7][14] ;
wire \d_pipe[7][15] ;
wire \d_pipe[7][16] ;
wire \d_pipe[7][17] ;
wire \d_pipe[7][18] ;
wire \d_pipe[7][19] ;
wire \d_pipe[7][20] ;
wire \d_pipe[7][21] ;
wire \d_pipe[7][22] ;
wire \d_pipe[7][23] ;
wire \d_pipe[8][12] ;
wire \d_pipe[8][13] ;
wire \d_pipe[8][14] ;
wire \d_pipe[8][15] ;
wire \d_pipe[8][16] ;
wire \d_pipe[8][17] ;
wire \d_pipe[8][18] ;
wire \d_pipe[8][19] ;
wire \d_pipe[8][20] ;
wire \d_pipe[8][21] ;
wire \d_pipe[8][22] ;
wire \d_pipe[8][23] ;
wire \d_pipe[9][12] ;
wire \q_pipe[10][0] ;
wire \q_pipe[10][1] ;
wire \q_pipe[10][2] ;
wire \q_pipe[10][3] ;
wire \q_pipe[10][4] ;
wire \q_pipe[10][5] ;
wire \q_pipe[10][6] ;
wire \q_pipe[10][7] ;
wire \q_pipe[10][8] ;
wire \q_pipe[10][9] ;
wire \q_pipe[11][0] ;
wire \q_pipe[11][10] ;
wire \q_pipe[11][1] ;
wire \q_pipe[11][2] ;
wire \q_pipe[11][3] ;
wire \q_pipe[11][4] ;
wire \q_pipe[11][5] ;
wire \q_pipe[11][6] ;
wire \q_pipe[11][7] ;
wire \q_pipe[11][8] ;
wire \q_pipe[11][9] ;
wire \q_pipe[1] ;
wire \q_pipe[2][0] ;
wire \q_pipe[2][1] ;
wire \q_pipe[3][0] ;
wire \q_pipe[3][1] ;
wire \q_pipe[3][2] ;
wire \q_pipe[4][0] ;
wire \q_pipe[4][1] ;
wire \q_pipe[4][2] ;
wire \q_pipe[4][3] ;
wire \q_pipe[5][0] ;
wire \q_pipe[5][1] ;
wire \q_pipe[5][2] ;
wire \q_pipe[5][3] ;
wire \q_pipe[5][4] ;
wire \q_pipe[6][0] ;
wire \q_pipe[6][1] ;
wire \q_pipe[6][2] ;
wire \q_pipe[6][3] ;
wire \q_pipe[6][4] ;
wire \q_pipe[6][5] ;
wire \q_pipe[7][0] ;
wire \q_pipe[7][1] ;
wire \q_pipe[7][2] ;
wire \q_pipe[7][3] ;
wire \q_pipe[7][4] ;
wire \q_pipe[7][5] ;
wire \q_pipe[7][6] ;
wire \q_pipe[8][0] ;
wire \q_pipe[8][1] ;
wire \q_pipe[8][2] ;
wire \q_pipe[8][3] ;
wire \q_pipe[8][4] ;
wire \q_pipe[8][5] ;
wire \q_pipe[8][6] ;
wire \q_pipe[8][7] ;
wire \q_pipe[9] ;
wire \s_pipe[10][10] ;
wire \s_pipe[10][11] ;
wire \s_pipe[10][12] ;
wire \s_pipe[10][13] ;
wire \s_pipe[10][14] ;
wire \s_pipe[10][15] ;
wire \s_pipe[10][16] ;
wire \s_pipe[10][17] ;
wire \s_pipe[10][18] ;
wire \s_pipe[10][19] ;
wire \s_pipe[10][20] ;
wire \s_pipe[10][21] ;
wire \s_pipe[10][22] ;
wire \s_pipe[10][23] ;
wire \s_pipe[10][24] ;
wire \s_pipe[11][11] ;
wire \s_pipe[11][12] ;
wire \s_pipe[11][13] ;
wire \s_pipe[11][14] ;
wire \s_pipe[11][15] ;
wire \s_pipe[11][16] ;
wire \s_pipe[11][17] ;
wire \s_pipe[11][18] ;
wire \s_pipe[11][19] ;
wire \s_pipe[11][20] ;
wire \s_pipe[11][21] ;
wire \s_pipe[11][22] ;
wire \s_pipe[11][23] ;
wire \s_pipe[11][24] ;
wire \s_pipe[12][24] ;
wire \s_pipe[1][10] ;
wire \s_pipe[1][11] ;
wire \s_pipe[1][12] ;
wire \s_pipe[1][13] ;
wire \s_pipe[1][14] ;
wire \s_pipe[1][15] ;
wire \s_pipe[1][16] ;
wire \s_pipe[1][17] ;
wire \s_pipe[1][18] ;
wire \s_pipe[1][19] ;
wire \s_pipe[1][1] ;
wire \s_pipe[1][20] ;
wire \s_pipe[1][21] ;
wire \s_pipe[1][22] ;
wire \s_pipe[1][23] ;
wire \s_pipe[1][24] ;
wire \s_pipe[1][2] ;
wire \s_pipe[1][3] ;
wire \s_pipe[1][4] ;
wire \s_pipe[1][5] ;
wire \s_pipe[1][6] ;
wire \s_pipe[1][7] ;
wire \s_pipe[1][8] ;
wire \s_pipe[1][9] ;
wire \s_pipe[2][10] ;
wire \s_pipe[2][11] ;
wire \s_pipe[2][12] ;
wire \s_pipe[2][13] ;
wire \s_pipe[2][14] ;
wire \s_pipe[2][15] ;
wire \s_pipe[2][16] ;
wire \s_pipe[2][17] ;
wire \s_pipe[2][18] ;
wire \s_pipe[2][19] ;
wire \s_pipe[2][20] ;
wire \s_pipe[2][21] ;
wire \s_pipe[2][22] ;
wire \s_pipe[2][23] ;
wire \s_pipe[2][24] ;
wire \s_pipe[2][2] ;
wire \s_pipe[2][3] ;
wire \s_pipe[2][4] ;
wire \s_pipe[2][5] ;
wire \s_pipe[2][6] ;
wire \s_pipe[2][7] ;
wire \s_pipe[2][8] ;
wire \s_pipe[2][9] ;
wire \s_pipe[3][10] ;
wire \s_pipe[3][11] ;
wire \s_pipe[3][12] ;
wire \s_pipe[3][13] ;
wire \s_pipe[3][14] ;
wire \s_pipe[3][15] ;
wire \s_pipe[3][16] ;
wire \s_pipe[3][17] ;
wire \s_pipe[3][18] ;
wire \s_pipe[3][19] ;
wire \s_pipe[3][20] ;
wire \s_pipe[3][21] ;
wire \s_pipe[3][22] ;
wire \s_pipe[3][23] ;
wire \s_pipe[3][24] ;
wire \s_pipe[3][3] ;
wire \s_pipe[3][4] ;
wire \s_pipe[3][5] ;
wire \s_pipe[3][6] ;
wire \s_pipe[3][7] ;
wire \s_pipe[3][8] ;
wire \s_pipe[3][9] ;
wire \s_pipe[4][10] ;
wire \s_pipe[4][11] ;
wire \s_pipe[4][12] ;
wire \s_pipe[4][13] ;
wire \s_pipe[4][14] ;
wire \s_pipe[4][15] ;
wire \s_pipe[4][16] ;
wire \s_pipe[4][17] ;
wire \s_pipe[4][18] ;
wire \s_pipe[4][19] ;
wire \s_pipe[4][20] ;
wire \s_pipe[4][21] ;
wire \s_pipe[4][22] ;
wire \s_pipe[4][23] ;
wire \s_pipe[4][24] ;
wire \s_pipe[4][4] ;
wire \s_pipe[4][5] ;
wire \s_pipe[4][6] ;
wire \s_pipe[4][7] ;
wire \s_pipe[4][8] ;
wire \s_pipe[4][9] ;
wire \s_pipe[5][10] ;
wire \s_pipe[5][11] ;
wire \s_pipe[5][12] ;
wire \s_pipe[5][13] ;
wire \s_pipe[5][14] ;
wire \s_pipe[5][15] ;
wire \s_pipe[5][16] ;
wire \s_pipe[5][17] ;
wire \s_pipe[5][18] ;
wire \s_pipe[5][19] ;
wire \s_pipe[5][20] ;
wire \s_pipe[5][21] ;
wire \s_pipe[5][22] ;
wire \s_pipe[5][23] ;
wire \s_pipe[5][24] ;
wire \s_pipe[5][5] ;
wire \s_pipe[5][6] ;
wire \s_pipe[5][7] ;
wire \s_pipe[5][8] ;
wire \s_pipe[5][9] ;
wire \s_pipe[6][10] ;
wire \s_pipe[6][11] ;
wire \s_pipe[6][12] ;
wire \s_pipe[6][13] ;
wire \s_pipe[6][14] ;
wire \s_pipe[6][15] ;
wire \s_pipe[6][16] ;
wire \s_pipe[6][17] ;
wire \s_pipe[6][18] ;
wire \s_pipe[6][19] ;
wire \s_pipe[6][20] ;
wire \s_pipe[6][21] ;
wire \s_pipe[6][22] ;
wire \s_pipe[6][23] ;
wire \s_pipe[6][24] ;
wire \s_pipe[6][6] ;
wire \s_pipe[6][7] ;
wire \s_pipe[6][8] ;
wire \s_pipe[6][9] ;
wire \s_pipe[7][10] ;
wire \s_pipe[7][11] ;
wire \s_pipe[7][12] ;
wire \s_pipe[7][13] ;
wire \s_pipe[7][14] ;
wire \s_pipe[7][15] ;
wire \s_pipe[7][16] ;
wire \s_pipe[7][17] ;
wire \s_pipe[7][18] ;
wire \s_pipe[7][19] ;
wire \s_pipe[7][20] ;
wire \s_pipe[7][21] ;
wire \s_pipe[7][22] ;
wire \s_pipe[7][23] ;
wire \s_pipe[7][24] ;
wire \s_pipe[7][7] ;
wire \s_pipe[7][8] ;
wire \s_pipe[7][9] ;
wire \s_pipe[8][10] ;
wire \s_pipe[8][11] ;
wire \s_pipe[8][12] ;
wire \s_pipe[8][13] ;
wire \s_pipe[8][14] ;
wire \s_pipe[8][15] ;
wire \s_pipe[8][16] ;
wire \s_pipe[8][17] ;
wire \s_pipe[8][18] ;
wire \s_pipe[8][19] ;
wire \s_pipe[8][20] ;
wire \s_pipe[8][21] ;
wire \s_pipe[8][22] ;
wire \s_pipe[8][23] ;
wire \s_pipe[8][24] ;
wire \s_pipe[8][8] ;
wire \s_pipe[8][9] ;
wire \s_pipe[9][10] ;
wire \s_pipe[9][11] ;
wire \s_pipe[9][12] ;
wire \s_pipe[9][13] ;
wire \s_pipe[9][14] ;
wire \s_pipe[9][9] ;

INV_X1 _4596_ (
  .A(\s_pipe[2][24] ),
  .ZN(_0626_)
);

NAND2_X1 _4597_ (
  .A1(_0626_),
  .A2(_4147_),
  .ZN(_0627_)
);

BUF_X2 _4598_ (
  .A(_0626_),
  .Z(_0628_)
);

OAI21_X1 _4599_ (
  .A(_0627_),
  .B1(_4145_),
  .B2(_0628_),
  .ZN(_4048_)
);

INV_X1 _4600_ (
  .A(_4048_),
  .ZN(_4044_)
);

INV_X1 _4601_ (
  .A(\s_pipe[3][24] ),
  .ZN(_0629_)
);

NAND2_X1 _4602_ (
  .A1(_0629_),
  .A2(_4183_),
  .ZN(_0630_)
);

BUF_X2 _4603_ (
  .A(_0629_),
  .Z(_0631_)
);

OAI21_X1 _4604_ (
  .A(_0630_),
  .B1(_4181_),
  .B2(_0631_),
  .ZN(_4055_)
);

INV_X1 _4605_ (
  .A(_4055_),
  .ZN(_4051_)
);

INV_X1 _4606_ (
  .A(\s_pipe[1][24] ),
  .ZN(_0632_)
);

BUF_X1 _4607_ (
  .A(_0632_),
  .Z(_0633_)
);

NAND2_X1 _4608_ (
  .A1(_0633_),
  .A2(_4219_),
  .ZN(_0634_)
);

OAI21_X1 _4609_ (
  .A(_0634_),
  .B1(_4217_),
  .B2(_0633_),
  .ZN(_4061_)
);

INV_X1 _4610_ (
  .A(_4061_),
  .ZN(_4057_)
);

INV_X1 _4611_ (
  .A(\s_pipe[11][24] ),
  .ZN(_0635_)
);

NAND2_X1 _4612_ (
  .A1(_0635_),
  .A2(_4288_),
  .ZN(_0636_)
);

BUF_X2 _4613_ (
  .A(_0635_),
  .Z(_0637_)
);

OAI21_X1 _4614_ (
  .A(_0636_),
  .B1(_4286_),
  .B2(_0637_),
  .ZN(_4071_)
);

INV_X1 _4615_ (
  .A(_4071_),
  .ZN(_4067_)
);

INV_X1 _4616_ (
  .A(\s_pipe[10][24] ),
  .ZN(_0638_)
);

BUF_X1 _4617_ (
  .A(_0638_),
  .Z(_0639_)
);

NAND2_X1 _4618_ (
  .A1(_0639_),
  .A2(_4324_),
  .ZN(_0640_)
);

OAI21_X1 _4619_ (
  .A(_0640_),
  .B1(_4322_),
  .B2(_0639_),
  .ZN(_4078_)
);

INV_X1 _4620_ (
  .A(_4078_),
  .ZN(_4074_)
);

BUF_X1 _4621_ (
  .A(_0000_),
  .Z(_0641_)
);

INV_X1 _4622_ (
  .A(_0641_),
  .ZN(_0642_)
);

BUF_X4 _4623_ (
  .A(_0642_),
  .Z(_0643_)
);

NAND2_X1 _4624_ (
  .A1(_0643_),
  .A2(_4360_),
  .ZN(_0644_)
);

OAI21_X1 _4625_ (
  .A(_0644_),
  .B1(_4358_),
  .B2(_0643_),
  .ZN(_4085_)
);

INV_X1 _4626_ (
  .A(_4085_),
  .ZN(_4081_)
);

INV_X1 _4627_ (
  .A(\s_pipe[8][24] ),
  .ZN(_0645_)
);

NAND2_X1 _4628_ (
  .A1(_0645_),
  .A2(_4396_),
  .ZN(_0646_)
);

BUF_X2 _4629_ (
  .A(_0645_),
  .Z(_0647_)
);

OAI21_X1 _4630_ (
  .A(_0646_),
  .B1(_4394_),
  .B2(_0647_),
  .ZN(_4092_)
);

INV_X1 _4631_ (
  .A(_4092_),
  .ZN(_4088_)
);

INV_X1 _4632_ (
  .A(\s_pipe[7][24] ),
  .ZN(_0648_)
);

NAND2_X1 _4633_ (
  .A1(_0648_),
  .A2(_4432_),
  .ZN(_0649_)
);

BUF_X1 _4634_ (
  .A(_0648_),
  .Z(_0650_)
);

OAI21_X1 _4635_ (
  .A(_0649_),
  .B1(_4430_),
  .B2(_0650_),
  .ZN(_4099_)
);

INV_X1 _4636_ (
  .A(_4099_),
  .ZN(_4095_)
);

INV_X1 _4637_ (
  .A(\s_pipe[6][24] ),
  .ZN(_0651_)
);

BUF_X2 _4638_ (
  .A(_0651_),
  .Z(_0652_)
);

NAND2_X1 _4639_ (
  .A1(_0652_),
  .A2(_4468_),
  .ZN(_0653_)
);

OAI21_X1 _4640_ (
  .A(_0653_),
  .B1(_4466_),
  .B2(_0652_),
  .ZN(_4106_)
);

INV_X1 _4641_ (
  .A(_4106_),
  .ZN(_4102_)
);

INV_X1 _4642_ (
  .A(\s_pipe[5][24] ),
  .ZN(_0654_)
);

BUF_X2 _4643_ (
  .A(_0654_),
  .Z(_0655_)
);

NAND2_X1 _4644_ (
  .A1(_0655_),
  .A2(_4504_),
  .ZN(_0656_)
);

OAI21_X1 _4645_ (
  .A(_0656_),
  .B1(_4502_),
  .B2(_0655_),
  .ZN(_4113_)
);

INV_X1 _4646_ (
  .A(_4113_),
  .ZN(_4109_)
);

INV_X1 _4647_ (
  .A(\s_pipe[4][24] ),
  .ZN(_0657_)
);

BUF_X2 _4648_ (
  .A(_0657_),
  .Z(_0658_)
);

NAND2_X1 _4649_ (
  .A1(_0658_),
  .A2(_4540_),
  .ZN(_0659_)
);

OAI21_X1 _4650_ (
  .A(_0659_),
  .B1(_4538_),
  .B2(_0658_),
  .ZN(_4120_)
);

INV_X1 _4651_ (
  .A(_4120_),
  .ZN(_4116_)
);

INV_X1 _4652_ (
  .A(z[12]),
  .ZN(_4063_)
);

INV_X1 _4653_ (
  .A(_4047_),
  .ZN(_4043_)
);

INV_X1 _4654_ (
  .A(_4054_),
  .ZN(_4050_)
);

INV_X1 _4655_ (
  .A(_4062_),
  .ZN(_4058_)
);

INV_X1 _4656_ (
  .A(_4072_),
  .ZN(_4068_)
);

INV_X1 _4657_ (
  .A(_4079_),
  .ZN(_4075_)
);

INV_X1 _4658_ (
  .A(_4086_),
  .ZN(_4082_)
);

INV_X1 _4659_ (
  .A(_4093_),
  .ZN(_4089_)
);

INV_X1 _4660_ (
  .A(_4100_),
  .ZN(_4096_)
);

INV_X1 _4661_ (
  .A(_4107_),
  .ZN(_4103_)
);

INV_X1 _4662_ (
  .A(_4114_),
  .ZN(_4110_)
);

INV_X1 _4663_ (
  .A(_4121_),
  .ZN(_4117_)
);

INV_X1 _4664_ (
  .A(z[11]),
  .ZN(_4122_)
);

INV_X1 _4665_ (
  .A(\d_pipe[2][13] ),
  .ZN(_0660_)
);

INV_X4 _4666_ (
  .A(\d_pipe[2][14] ),
  .ZN(_0661_)
);

AND3_X4 _4667_ (
  .A1(_0660_),
  .A2(_0661_),
  .A3(_4144_),
  .ZN(_0662_)
);

INV_X2 _4668_ (
  .A(\d_pipe[2][15] ),
  .ZN(_0663_)
);

OAI21_X1 _4669_ (
  .A(_0628_),
  .B1(_0662_),
  .B2(_0663_),
  .ZN(_0664_)
);

NAND2_X2 _4670_ (
  .A1(_0662_),
  .A2(_0663_),
  .ZN(_0665_)
);

INV_X1 _4671_ (
  .A(_0665_),
  .ZN(_0666_)
);

BUF_X1 _4672_ (
  .A(_0626_),
  .Z(_0667_)
);

OAI22_X1 _4673_ (
  .A1(_0664_),
  .A2(_0666_),
  .B1(_0092_),
  .B2(_0667_),
  .ZN(_4153_)
);

XNOR2_X1 _4674_ (
  .A(_4218_),
  .B(\d_pipe[1][14] ),
  .ZN(_0668_)
);

BUF_X1 _4675_ (
  .A(_0632_),
  .Z(_0669_)
);

NAND2_X1 _4676_ (
  .A1(_0668_),
  .A2(_0669_),
  .ZN(_0670_)
);

OAI21_X1 _4677_ (
  .A(_0670_),
  .B1(_0669_),
  .B2(_0001_),
  .ZN(_4222_)
);

INV_X2 _4678_ (
  .A(\d_pipe[1][14] ),
  .ZN(_0671_)
);

INV_X1 _4679_ (
  .A(\d_pipe[1][13] ),
  .ZN(_0672_)
);

NAND3_X1 _4680_ (
  .A1(_0671_),
  .A2(_0672_),
  .A3(_4216_),
  .ZN(_0673_)
);

INV_X1 _4681_ (
  .A(_0673_),
  .ZN(_0674_)
);

INV_X4 _4682_ (
  .A(\d_pipe[1][15] ),
  .ZN(_0675_)
);

OAI21_X1 _4683_ (
  .A(_0633_),
  .B1(_0674_),
  .B2(_0675_),
  .ZN(_0676_)
);

NAND2_X1 _4684_ (
  .A1(_0674_),
  .A2(_0675_),
  .ZN(_0677_)
);

INV_X1 _4685_ (
  .A(_0677_),
  .ZN(_0678_)
);

OAI22_X1 _4686_ (
  .A1(_0676_),
  .A2(_0678_),
  .B1(_0002_),
  .B2(_0669_),
  .ZN(_4225_)
);

INV_X2 _4687_ (
  .A(_3715_),
  .ZN(_0679_)
);

INV_X4 _4688_ (
  .A(_3716_),
  .ZN(_0680_)
);

NAND3_X2 _4689_ (
  .A1(_0679_),
  .A2(_0680_),
  .A3(_4359_),
  .ZN(_0681_)
);

BUF_X4 _4690_ (
  .A(_3717_),
  .Z(_0682_)
);

OR2_X1 _4691_ (
  .A1(_0681_),
  .A2(_0682_),
  .ZN(_0683_)
);

BUF_X4 _4692_ (
  .A(_0643_),
  .Z(_0684_)
);

NAND2_X1 _4693_ (
  .A1(_0681_),
  .A2(_0682_),
  .ZN(_0685_)
);

NAND3_X1 _4694_ (
  .A1(_0683_),
  .A2(_0684_),
  .A3(_0685_),
  .ZN(_0686_)
);

OAI21_X1 _4695_ (
  .A(_0686_),
  .B1(_0684_),
  .B2(_0033_),
  .ZN(_4369_)
);

XNOR2_X1 _4696_ (
  .A(_4146_),
  .B(\d_pipe[2][14] ),
  .ZN(_0687_)
);

NAND2_X1 _4697_ (
  .A1(_0687_),
  .A2(_0667_),
  .ZN(_0688_)
);

OAI21_X1 _4698_ (
  .A(_0688_),
  .B1(_0667_),
  .B2(_0091_),
  .ZN(_4150_)
);

NAND3_X4 _4699_ (
  .A1(_0661_),
  .A2(_0663_),
  .A3(_4146_),
  .ZN(_0689_)
);

BUF_X4 _4700_ (
  .A(\d_pipe[2][16] ),
  .Z(_0690_)
);

OR2_X1 _4701_ (
  .A1(_0689_),
  .A2(_0690_),
  .ZN(_0691_)
);

NAND2_X1 _4702_ (
  .A1(_0689_),
  .A2(_0690_),
  .ZN(_0692_)
);

NAND3_X1 _4703_ (
  .A1(_0691_),
  .A2(_0628_),
  .A3(_0692_),
  .ZN(_0693_)
);

OAI21_X1 _4704_ (
  .A(_0693_),
  .B1(_0667_),
  .B2(_0093_),
  .ZN(_4156_)
);

NOR2_X4 _4705_ (
  .A1(_0665_),
  .A2(_0690_),
  .ZN(_0694_)
);

BUF_X4 _4706_ (
  .A(\d_pipe[2][17] ),
  .Z(_0695_)
);

INV_X2 _4707_ (
  .A(_0695_),
  .ZN(_0696_)
);

NAND2_X2 _4708_ (
  .A1(_0694_),
  .A2(_0696_),
  .ZN(_0697_)
);

OAI21_X1 _4709_ (
  .A(_0695_),
  .B1(_0665_),
  .B2(_0690_),
  .ZN(_0698_)
);

NAND3_X1 _4710_ (
  .A1(_0697_),
  .A2(_0698_),
  .A3(_0628_),
  .ZN(_0699_)
);

OAI21_X1 _4711_ (
  .A(_0699_),
  .B1(_0667_),
  .B2(_0094_),
  .ZN(_4159_)
);

NOR2_X1 _4712_ (
  .A1(_0691_),
  .A2(_0695_),
  .ZN(_0700_)
);

BUF_X4 _4713_ (
  .A(\d_pipe[2][18] ),
  .Z(_0701_)
);

INV_X2 _4714_ (
  .A(_0701_),
  .ZN(_0702_)
);

OAI21_X1 _4715_ (
  .A(_0628_),
  .B1(_0700_),
  .B2(_0702_),
  .ZN(_0703_)
);

NOR3_X1 _4716_ (
  .A1(_0691_),
  .A2(_0695_),
  .A3(_0701_),
  .ZN(_0704_)
);

OAI22_X1 _4717_ (
  .A1(_0703_),
  .A2(_0704_),
  .B1(_0095_),
  .B2(_0667_),
  .ZN(_4162_)
);

NOR2_X1 _4718_ (
  .A1(_0697_),
  .A2(_0701_),
  .ZN(_0705_)
);

INV_X1 _4719_ (
  .A(\d_pipe[2][19] ),
  .ZN(_0706_)
);

NOR2_X1 _4720_ (
  .A1(_0705_),
  .A2(_0706_),
  .ZN(_0707_)
);

NOR2_X4 _4721_ (
  .A1(_0701_),
  .A2(\d_pipe[2][19] ),
  .ZN(_0708_)
);

NAND3_X1 _4722_ (
  .A1(_0694_),
  .A2(_0696_),
  .A3(_0708_),
  .ZN(_0709_)
);

NAND2_X1 _4723_ (
  .A1(_0709_),
  .A2(_0628_),
  .ZN(_0710_)
);

OAI22_X1 _4724_ (
  .A1(_0707_),
  .A2(_0710_),
  .B1(_0096_),
  .B2(_0667_),
  .ZN(_4165_)
);

OR2_X1 _4725_ (
  .A1(_0628_),
  .A2(_0097_),
  .ZN(_0711_)
);

NOR2_X4 _4726_ (
  .A1(_0690_),
  .A2(_0695_),
  .ZN(_0712_)
);

NAND2_X2 _4727_ (
  .A1(_0712_),
  .A2(_0708_),
  .ZN(_0713_)
);

NOR2_X4 _4728_ (
  .A1(_0713_),
  .A2(_0689_),
  .ZN(_0714_)
);

INV_X1 _4729_ (
  .A(\d_pipe[2][20] ),
  .ZN(_0715_)
);

XNOR2_X1 _4730_ (
  .A(_0714_),
  .B(_0715_),
  .ZN(_0716_)
);

OAI21_X1 _4731_ (
  .A(_0711_),
  .B1(_0716_),
  .B2(\s_pipe[2][24] ),
  .ZN(_4168_)
);

INV_X2 _4732_ (
  .A(_0690_),
  .ZN(_0717_)
);

NAND4_X1 _4733_ (
  .A1(_0663_),
  .A2(_0717_),
  .A3(_0661_),
  .A4(_0660_),
  .ZN(_0718_)
);

NAND2_X1 _4734_ (
  .A1(_0696_),
  .A2(_0702_),
  .ZN(_0719_)
);

NAND2_X1 _4735_ (
  .A1(_0706_),
  .A2(_0715_),
  .ZN(_0720_)
);

NOR3_X2 _4736_ (
  .A1(_0718_),
  .A2(_0719_),
  .A3(_0720_),
  .ZN(_0721_)
);

BUF_X4 _4737_ (
  .A(\d_pipe[2][21] ),
  .Z(_0722_)
);

NAND3_X1 _4738_ (
  .A1(_0721_),
  .A2(_4144_),
  .A3(_0722_),
  .ZN(_0723_)
);

INV_X1 _4739_ (
  .A(_0723_),
  .ZN(_0724_)
);

AOI21_X1 _4740_ (
  .A(_0722_),
  .B1(_0721_),
  .B2(_4144_),
  .ZN(_0725_)
);

OAI21_X1 _4741_ (
  .A(_0667_),
  .B1(_0724_),
  .B2(_0725_),
  .ZN(_0726_)
);

OR2_X1 _4742_ (
  .A1(_0628_),
  .A2(_0098_),
  .ZN(_0727_)
);

NAND2_X1 _4743_ (
  .A1(_0726_),
  .A2(_0727_),
  .ZN(_4171_)
);

INV_X1 _4744_ (
  .A(_0714_),
  .ZN(_0728_)
);

NOR2_X4 _4745_ (
  .A1(\d_pipe[2][20] ),
  .A2(_0722_),
  .ZN(_0729_)
);

INV_X1 _4746_ (
  .A(\d_pipe[2][22] ),
  .ZN(_0730_)
);

NAND2_X2 _4747_ (
  .A1(_0729_),
  .A2(_0730_),
  .ZN(_0731_)
);

OAI21_X1 _4748_ (
  .A(_0628_),
  .B1(_0728_),
  .B2(_0731_),
  .ZN(_0732_)
);

AOI21_X1 _4749_ (
  .A(_0730_),
  .B1(_0714_),
  .B2(_0729_),
  .ZN(_0733_)
);

OAI22_X1 _4750_ (
  .A1(_0732_),
  .A2(_0733_),
  .B1(_0099_),
  .B2(_0667_),
  .ZN(_4174_)
);

NAND4_X1 _4751_ (
  .A1(_0696_),
  .A2(_0702_),
  .A3(_0663_),
  .A4(_0717_),
  .ZN(_0734_)
);

INV_X1 _4752_ (
  .A(_0722_),
  .ZN(_0735_)
);

NAND2_X1 _4753_ (
  .A1(_0735_),
  .A2(_0730_),
  .ZN(_0736_)
);

NOR3_X2 _4754_ (
  .A1(_0734_),
  .A2(_0720_),
  .A3(_0736_),
  .ZN(_0737_)
);

BUF_X1 _4755_ (
  .A(\d_pipe[2][23] ),
  .Z(_0738_)
);

NAND3_X1 _4756_ (
  .A1(_0737_),
  .A2(_0738_),
  .A3(_0662_),
  .ZN(_0739_)
);

INV_X1 _4757_ (
  .A(_0739_),
  .ZN(_0740_)
);

AOI21_X1 _4758_ (
  .A(_0738_),
  .B1(_0737_),
  .B2(_0662_),
  .ZN(_0741_)
);

OAI21_X1 _4759_ (
  .A(_0667_),
  .B1(_0740_),
  .B2(_0741_),
  .ZN(_0742_)
);

OR2_X1 _4760_ (
  .A1(_0628_),
  .A2(_0100_),
  .ZN(_0743_)
);

NAND2_X1 _4761_ (
  .A1(_0742_),
  .A2(_0743_),
  .ZN(_4177_)
);

XNOR2_X1 _4762_ (
  .A(_4182_),
  .B(\d_pipe[3][14] ),
  .ZN(_0744_)
);

BUF_X1 _4763_ (
  .A(_0629_),
  .Z(_0745_)
);

NAND2_X1 _4764_ (
  .A1(_0744_),
  .A2(_0745_),
  .ZN(_0746_)
);

OAI21_X1 _4765_ (
  .A(_0746_),
  .B1(_0745_),
  .B2(_0101_),
  .ZN(_4186_)
);

INV_X4 _4766_ (
  .A(\d_pipe[3][14] ),
  .ZN(_0747_)
);

INV_X2 _4767_ (
  .A(\d_pipe[3][13] ),
  .ZN(_0748_)
);

NAND3_X2 _4768_ (
  .A1(_0747_),
  .A2(_0748_),
  .A3(_4180_),
  .ZN(_0749_)
);

INV_X2 _4769_ (
  .A(_0749_),
  .ZN(_0750_)
);

INV_X4 _4770_ (
  .A(\d_pipe[3][15] ),
  .ZN(_0751_)
);

OAI21_X1 _4771_ (
  .A(_0631_),
  .B1(_0750_),
  .B2(_0751_),
  .ZN(_0752_)
);

NAND2_X1 _4772_ (
  .A1(_0750_),
  .A2(_0751_),
  .ZN(_0753_)
);

INV_X1 _4773_ (
  .A(_0753_),
  .ZN(_0754_)
);

OAI22_X1 _4774_ (
  .A1(_0752_),
  .A2(_0754_),
  .B1(_0102_),
  .B2(_0745_),
  .ZN(_4189_)
);

NAND3_X2 _4775_ (
  .A1(_0747_),
  .A2(_0751_),
  .A3(_4182_),
  .ZN(_0755_)
);

BUF_X2 _4776_ (
  .A(\d_pipe[3][16] ),
  .Z(_0756_)
);

OR2_X1 _4777_ (
  .A1(_0755_),
  .A2(_0756_),
  .ZN(_0757_)
);

NAND2_X1 _4778_ (
  .A1(_0755_),
  .A2(_0756_),
  .ZN(_0758_)
);

NAND3_X1 _4779_ (
  .A1(_0757_),
  .A2(_0631_),
  .A3(_0758_),
  .ZN(_0759_)
);

OAI21_X1 _4780_ (
  .A(_0759_),
  .B1(_0745_),
  .B2(_0103_),
  .ZN(_4192_)
);

INV_X2 _4781_ (
  .A(_0756_),
  .ZN(_0760_)
);

NAND2_X1 _4782_ (
  .A1(_0754_),
  .A2(_0760_),
  .ZN(_0761_)
);

INV_X1 _4783_ (
  .A(_0761_),
  .ZN(_0762_)
);

BUF_X4 _4784_ (
  .A(\d_pipe[3][17] ),
  .Z(_0763_)
);

INV_X1 _4785_ (
  .A(_0763_),
  .ZN(_0764_)
);

OAI21_X1 _4786_ (
  .A(_0631_),
  .B1(_0762_),
  .B2(_0764_),
  .ZN(_0765_)
);

NOR2_X2 _4787_ (
  .A1(_0761_),
  .A2(_0763_),
  .ZN(_0766_)
);

OAI22_X1 _4788_ (
  .A1(_0765_),
  .A2(_0766_),
  .B1(_0104_),
  .B2(_0745_),
  .ZN(_4195_)
);

NOR2_X1 _4789_ (
  .A1(_0757_),
  .A2(_0763_),
  .ZN(_0767_)
);

INV_X1 _4790_ (
  .A(\d_pipe[3][18] ),
  .ZN(_0768_)
);

OAI21_X1 _4791_ (
  .A(_0631_),
  .B1(_0767_),
  .B2(_0768_),
  .ZN(_0769_)
);

NOR3_X1 _4792_ (
  .A1(_0757_),
  .A2(_0763_),
  .A3(\d_pipe[3][18] ),
  .ZN(_0770_)
);

OAI22_X1 _4793_ (
  .A1(_0769_),
  .A2(_0770_),
  .B1(_0105_),
  .B2(_0745_),
  .ZN(_4198_)
);

NOR2_X2 _4794_ (
  .A1(\d_pipe[3][18] ),
  .A2(\d_pipe[3][19] ),
  .ZN(_0771_)
);

NAND2_X1 _4795_ (
  .A1(_0766_),
  .A2(_0771_),
  .ZN(_0772_)
);

NAND4_X2 _4796_ (
  .A1(_0764_),
  .A2(_0768_),
  .A3(_0751_),
  .A4(_0760_),
  .ZN(_0773_)
);

OAI21_X1 _4797_ (
  .A(\d_pipe[3][19] ),
  .B1(_0773_),
  .B2(_0749_),
  .ZN(_0774_)
);

NAND3_X1 _4798_ (
  .A1(_0772_),
  .A2(_0631_),
  .A3(_0774_),
  .ZN(_0775_)
);

OAI21_X1 _4799_ (
  .A(_0775_),
  .B1(_0745_),
  .B2(_0106_),
  .ZN(_4201_)
);

OR2_X1 _4800_ (
  .A1(_0631_),
  .A2(_0107_),
  .ZN(_0776_)
);

NOR2_X4 _4801_ (
  .A1(_0756_),
  .A2(_0763_),
  .ZN(_0777_)
);

NAND2_X2 _4802_ (
  .A1(_0777_),
  .A2(_0771_),
  .ZN(_0778_)
);

NOR2_X4 _4803_ (
  .A1(_0778_),
  .A2(_0755_),
  .ZN(_0779_)
);

INV_X1 _4804_ (
  .A(\d_pipe[3][20] ),
  .ZN(_0780_)
);

XNOR2_X1 _4805_ (
  .A(_0779_),
  .B(_0780_),
  .ZN(_0781_)
);

OAI21_X1 _4806_ (
  .A(_0776_),
  .B1(_0781_),
  .B2(\s_pipe[3][24] ),
  .ZN(_4204_)
);

NAND4_X1 _4807_ (
  .A1(_0751_),
  .A2(_0760_),
  .A3(_0747_),
  .A4(_0748_),
  .ZN(_0782_)
);

NAND2_X1 _4808_ (
  .A1(_0764_),
  .A2(_0768_),
  .ZN(_0783_)
);

INV_X1 _4809_ (
  .A(\d_pipe[3][19] ),
  .ZN(_0784_)
);

NAND2_X1 _4810_ (
  .A1(_0784_),
  .A2(_0780_),
  .ZN(_0785_)
);

NOR3_X2 _4811_ (
  .A1(_0782_),
  .A2(_0783_),
  .A3(_0785_),
  .ZN(_0786_)
);

NAND2_X1 _4812_ (
  .A1(_0786_),
  .A2(_4180_),
  .ZN(_0787_)
);

NAND2_X1 _4813_ (
  .A1(_0787_),
  .A2(\d_pipe[3][21] ),
  .ZN(_0788_)
);

INV_X1 _4814_ (
  .A(\d_pipe[3][21] ),
  .ZN(_0789_)
);

NAND3_X1 _4815_ (
  .A1(_0786_),
  .A2(_4180_),
  .A3(_0789_),
  .ZN(_0790_)
);

NAND3_X1 _4816_ (
  .A1(_0788_),
  .A2(_0790_),
  .A3(_0631_),
  .ZN(_0791_)
);

OAI21_X1 _4817_ (
  .A(_0791_),
  .B1(_0745_),
  .B2(_0108_),
  .ZN(_4207_)
);

INV_X1 _4818_ (
  .A(_0779_),
  .ZN(_0792_)
);

NOR2_X2 _4819_ (
  .A1(\d_pipe[3][20] ),
  .A2(\d_pipe[3][21] ),
  .ZN(_0793_)
);

INV_X1 _4820_ (
  .A(\d_pipe[3][22] ),
  .ZN(_0794_)
);

NAND2_X1 _4821_ (
  .A1(_0793_),
  .A2(_0794_),
  .ZN(_0795_)
);

OAI21_X1 _4822_ (
  .A(_0631_),
  .B1(_0792_),
  .B2(_0795_),
  .ZN(_0796_)
);

AOI21_X1 _4823_ (
  .A(_0794_),
  .B1(_0779_),
  .B2(_0793_),
  .ZN(_0797_)
);

OAI22_X1 _4824_ (
  .A1(_0796_),
  .A2(_0797_),
  .B1(_0109_),
  .B2(_0745_),
  .ZN(_4210_)
);

NAND4_X1 _4825_ (
  .A1(_0789_),
  .A2(_0794_),
  .A3(_0784_),
  .A4(_0780_),
  .ZN(_0798_)
);

NOR2_X2 _4826_ (
  .A1(_0773_),
  .A2(_0798_),
  .ZN(_0799_)
);

INV_X1 _4827_ (
  .A(_0799_),
  .ZN(_0800_)
);

OAI21_X1 _4828_ (
  .A(\d_pipe[3][23] ),
  .B1(_0800_),
  .B2(_0749_),
  .ZN(_0801_)
);

INV_X1 _4829_ (
  .A(\d_pipe[3][23] ),
  .ZN(_0802_)
);

NAND3_X1 _4830_ (
  .A1(_0799_),
  .A2(_0802_),
  .A3(_0750_),
  .ZN(_0803_)
);

NAND3_X1 _4831_ (
  .A1(_0801_),
  .A2(_0631_),
  .A3(_0803_),
  .ZN(_0804_)
);

OAI21_X1 _4832_ (
  .A(_0804_),
  .B1(_0745_),
  .B2(_0110_),
  .ZN(_4213_)
);

NAND3_X2 _4833_ (
  .A1(_0671_),
  .A2(_0675_),
  .A3(_4218_),
  .ZN(_0805_)
);

BUF_X4 _4834_ (
  .A(\d_pipe[1][16] ),
  .Z(_0806_)
);

OR2_X1 _4835_ (
  .A1(_0805_),
  .A2(_0806_),
  .ZN(_0807_)
);

NAND2_X1 _4836_ (
  .A1(_0805_),
  .A2(_0806_),
  .ZN(_0808_)
);

NAND3_X1 _4837_ (
  .A1(_0807_),
  .A2(_0633_),
  .A3(_0808_),
  .ZN(_0809_)
);

OAI21_X1 _4838_ (
  .A(_0809_),
  .B1(_0669_),
  .B2(_0003_),
  .ZN(_4228_)
);

INV_X2 _4839_ (
  .A(_0806_),
  .ZN(_0810_)
);

BUF_X4 _4840_ (
  .A(\d_pipe[1][17] ),
  .Z(_0811_)
);

INV_X2 _4841_ (
  .A(_0811_),
  .ZN(_0812_)
);

NAND3_X1 _4842_ (
  .A1(_0678_),
  .A2(_0810_),
  .A3(_0812_),
  .ZN(_0813_)
);

OAI21_X1 _4843_ (
  .A(_0811_),
  .B1(_0677_),
  .B2(_0806_),
  .ZN(_0814_)
);

NAND3_X1 _4844_ (
  .A1(_0813_),
  .A2(_0814_),
  .A3(_0633_),
  .ZN(_0815_)
);

OAI21_X1 _4845_ (
  .A(_0815_),
  .B1(_0669_),
  .B2(_0004_),
  .ZN(_4231_)
);

NOR2_X1 _4846_ (
  .A1(_0807_),
  .A2(_0811_),
  .ZN(_0816_)
);

INV_X1 _4847_ (
  .A(\d_pipe[1][18] ),
  .ZN(_0817_)
);

OAI21_X1 _4848_ (
  .A(_0633_),
  .B1(_0816_),
  .B2(_0817_),
  .ZN(_0818_)
);

NOR3_X1 _4849_ (
  .A1(_0807_),
  .A2(_0811_),
  .A3(\d_pipe[1][18] ),
  .ZN(_0819_)
);

OAI22_X1 _4850_ (
  .A1(_0818_),
  .A2(_0819_),
  .B1(_0005_),
  .B2(_0669_),
  .ZN(_4234_)
);

OR2_X1 _4851_ (
  .A1(_0633_),
  .A2(_0006_),
  .ZN(_0820_)
);

NAND4_X2 _4852_ (
  .A1(_0812_),
  .A2(_0817_),
  .A3(_0675_),
  .A4(_0810_),
  .ZN(_0821_)
);

NOR2_X1 _4853_ (
  .A1(_0821_),
  .A2(_0673_),
  .ZN(_0822_)
);

INV_X1 _4854_ (
  .A(\d_pipe[1][19] ),
  .ZN(_0823_)
);

XNOR2_X1 _4855_ (
  .A(_0822_),
  .B(_0823_),
  .ZN(_0824_)
);

OAI21_X1 _4856_ (
  .A(_0820_),
  .B1(_0824_),
  .B2(\s_pipe[1][24] ),
  .ZN(_4237_)
);

OR2_X1 _4857_ (
  .A1(_0633_),
  .A2(_0007_),
  .ZN(_0825_)
);

NOR2_X4 _4858_ (
  .A1(_0806_),
  .A2(_0811_),
  .ZN(_0826_)
);

NOR2_X1 _4859_ (
  .A1(\d_pipe[1][18] ),
  .A2(\d_pipe[1][19] ),
  .ZN(_0827_)
);

NAND2_X2 _4860_ (
  .A1(_0826_),
  .A2(_0827_),
  .ZN(_0828_)
);

NOR2_X4 _4861_ (
  .A1(_0828_),
  .A2(_0805_),
  .ZN(_0829_)
);

INV_X1 _4862_ (
  .A(\d_pipe[1][20] ),
  .ZN(_0830_)
);

XNOR2_X1 _4863_ (
  .A(_0829_),
  .B(_0830_),
  .ZN(_0831_)
);

OAI21_X1 _4864_ (
  .A(_0825_),
  .B1(_0831_),
  .B2(\s_pipe[1][24] ),
  .ZN(_4240_)
);

NAND4_X1 _4865_ (
  .A1(_0675_),
  .A2(_0810_),
  .A3(_0671_),
  .A4(_0672_),
  .ZN(_0832_)
);

NAND2_X1 _4866_ (
  .A1(_0812_),
  .A2(_0817_),
  .ZN(_0833_)
);

NAND2_X1 _4867_ (
  .A1(_0823_),
  .A2(_0830_),
  .ZN(_0834_)
);

NOR3_X2 _4868_ (
  .A1(_0832_),
  .A2(_0833_),
  .A3(_0834_),
  .ZN(_0835_)
);

NAND2_X1 _4869_ (
  .A1(_0835_),
  .A2(_4216_),
  .ZN(_0836_)
);

NAND2_X1 _4870_ (
  .A1(_0836_),
  .A2(\d_pipe[1][21] ),
  .ZN(_0837_)
);

INV_X1 _4871_ (
  .A(\d_pipe[1][21] ),
  .ZN(_0838_)
);

NAND3_X1 _4872_ (
  .A1(_0835_),
  .A2(_4216_),
  .A3(_0838_),
  .ZN(_0839_)
);

NAND3_X1 _4873_ (
  .A1(_0837_),
  .A2(_0839_),
  .A3(_0633_),
  .ZN(_0840_)
);

OAI21_X1 _4874_ (
  .A(_0840_),
  .B1(_0669_),
  .B2(_0008_),
  .ZN(_4243_)
);

INV_X1 _4875_ (
  .A(_0829_),
  .ZN(_0841_)
);

NOR2_X2 _4876_ (
  .A1(\d_pipe[1][20] ),
  .A2(\d_pipe[1][21] ),
  .ZN(_0842_)
);

INV_X1 _4877_ (
  .A(\d_pipe[1][22] ),
  .ZN(_0843_)
);

NAND2_X1 _4878_ (
  .A1(_0842_),
  .A2(_0843_),
  .ZN(_0844_)
);

OAI21_X1 _4879_ (
  .A(_0633_),
  .B1(_0841_),
  .B2(_0844_),
  .ZN(_0845_)
);

AOI21_X1 _4880_ (
  .A(_0843_),
  .B1(_0829_),
  .B2(_0842_),
  .ZN(_0846_)
);

OAI22_X1 _4881_ (
  .A1(_0845_),
  .A2(_0846_),
  .B1(_0009_),
  .B2(_0669_),
  .ZN(_4246_)
);

NAND4_X1 _4882_ (
  .A1(_0838_),
  .A2(_0843_),
  .A3(_0823_),
  .A4(_0830_),
  .ZN(_0847_)
);

NOR2_X2 _4883_ (
  .A1(_0821_),
  .A2(_0847_),
  .ZN(_0848_)
);

INV_X1 _4884_ (
  .A(_0848_),
  .ZN(_0849_)
);

OAI21_X1 _4885_ (
  .A(\d_pipe[1][23] ),
  .B1(_0849_),
  .B2(_0673_),
  .ZN(_0850_)
);

INV_X1 _4886_ (
  .A(\d_pipe[1][23] ),
  .ZN(_0851_)
);

NAND3_X1 _4887_ (
  .A1(_0848_),
  .A2(_0851_),
  .A3(_0674_),
  .ZN(_0852_)
);

NAND3_X1 _4888_ (
  .A1(_0850_),
  .A2(_0669_),
  .A3(_0852_),
  .ZN(_0853_)
);

OAI21_X1 _4889_ (
  .A(_0853_),
  .B1(_0669_),
  .B2(_0010_),
  .ZN(_4249_)
);

INV_X1 _4890_ (
  .A(d[2]),
  .ZN(_4255_)
);

INV_X1 _4891_ (
  .A(d[5]),
  .ZN(_4264_)
);

INV_X1 _4892_ (
  .A(d[6]),
  .ZN(_4267_)
);

INV_X1 _4893_ (
  .A(d[7]),
  .ZN(_4270_)
);

INV_X1 _4894_ (
  .A(d[8]),
  .ZN(_4273_)
);

INV_X1 _4895_ (
  .A(d[9]),
  .ZN(_4276_)
);

XNOR2_X1 _4896_ (
  .A(_4287_),
  .B(\d_pipe[11][14] ),
  .ZN(_0854_)
);

BUF_X1 _4897_ (
  .A(_0635_),
  .Z(_0855_)
);

NAND2_X1 _4898_ (
  .A1(_0854_),
  .A2(_0855_),
  .ZN(_0856_)
);

OAI21_X1 _4899_ (
  .A(_0856_),
  .B1(_0855_),
  .B2(_0011_),
  .ZN(_4291_)
);

INV_X2 _4900_ (
  .A(\d_pipe[11][14] ),
  .ZN(_0857_)
);

INV_X2 _4901_ (
  .A(\d_pipe[11][13] ),
  .ZN(_0858_)
);

NAND3_X2 _4902_ (
  .A1(_0857_),
  .A2(_0858_),
  .A3(_4285_),
  .ZN(_0859_)
);

INV_X2 _4903_ (
  .A(_0859_),
  .ZN(_0860_)
);

INV_X4 _4904_ (
  .A(\d_pipe[11][15] ),
  .ZN(_0861_)
);

OAI21_X1 _4905_ (
  .A(_0637_),
  .B1(_0860_),
  .B2(_0861_),
  .ZN(_0862_)
);

NAND2_X1 _4906_ (
  .A1(_0860_),
  .A2(_0861_),
  .ZN(_0863_)
);

INV_X1 _4907_ (
  .A(_0863_),
  .ZN(_0864_)
);

OAI22_X1 _4908_ (
  .A1(_0862_),
  .A2(_0864_),
  .B1(_0012_),
  .B2(_0855_),
  .ZN(_4294_)
);

NAND3_X2 _4909_ (
  .A1(_0857_),
  .A2(_0861_),
  .A3(_4287_),
  .ZN(_0865_)
);

OR2_X1 _4910_ (
  .A1(_0865_),
  .A2(\d_pipe[11][16] ),
  .ZN(_0866_)
);

NAND2_X1 _4911_ (
  .A1(_0865_),
  .A2(\d_pipe[11][16] ),
  .ZN(_0867_)
);

NAND3_X1 _4912_ (
  .A1(_0866_),
  .A2(_0637_),
  .A3(_0867_),
  .ZN(_0868_)
);

OAI21_X1 _4913_ (
  .A(_0868_),
  .B1(_0855_),
  .B2(_0013_),
  .ZN(_4297_)
);

INV_X2 _4914_ (
  .A(\d_pipe[11][16] ),
  .ZN(_0869_)
);

NAND2_X1 _4915_ (
  .A1(_0864_),
  .A2(_0869_),
  .ZN(_0870_)
);

INV_X1 _4916_ (
  .A(_0870_),
  .ZN(_0871_)
);

BUF_X4 _4917_ (
  .A(\d_pipe[11][17] ),
  .Z(_0872_)
);

INV_X2 _4918_ (
  .A(_0872_),
  .ZN(_0873_)
);

OAI21_X1 _4919_ (
  .A(_0637_),
  .B1(_0871_),
  .B2(_0873_),
  .ZN(_0874_)
);

NOR2_X2 _4920_ (
  .A1(_0870_),
  .A2(_0872_),
  .ZN(_0875_)
);

OAI22_X1 _4921_ (
  .A1(_0874_),
  .A2(_0875_),
  .B1(_0014_),
  .B2(_0855_),
  .ZN(_4300_)
);

NOR2_X1 _4922_ (
  .A1(_0866_),
  .A2(_0872_),
  .ZN(_0876_)
);

INV_X1 _4923_ (
  .A(\d_pipe[11][18] ),
  .ZN(_0877_)
);

OAI21_X1 _4924_ (
  .A(_0637_),
  .B1(_0876_),
  .B2(_0877_),
  .ZN(_0878_)
);

NOR3_X1 _4925_ (
  .A1(_0866_),
  .A2(_0872_),
  .A3(\d_pipe[11][18] ),
  .ZN(_0879_)
);

OAI22_X1 _4926_ (
  .A1(_0878_),
  .A2(_0879_),
  .B1(_0015_),
  .B2(_0855_),
  .ZN(_4303_)
);

NOR2_X2 _4927_ (
  .A1(\d_pipe[11][18] ),
  .A2(\d_pipe[11][19] ),
  .ZN(_0880_)
);

NAND2_X1 _4928_ (
  .A1(_0875_),
  .A2(_0880_),
  .ZN(_0881_)
);

NAND4_X1 _4929_ (
  .A1(_0873_),
  .A2(_0877_),
  .A3(_0861_),
  .A4(_0869_),
  .ZN(_0882_)
);

OAI21_X1 _4930_ (
  .A(\d_pipe[11][19] ),
  .B1(_0882_),
  .B2(_0859_),
  .ZN(_0883_)
);

NAND3_X1 _4931_ (
  .A1(_0881_),
  .A2(_0637_),
  .A3(_0883_),
  .ZN(_0884_)
);

OAI21_X1 _4932_ (
  .A(_0884_),
  .B1(_0855_),
  .B2(_0016_),
  .ZN(_4306_)
);

OR2_X1 _4933_ (
  .A1(_0637_),
  .A2(_0017_),
  .ZN(_0885_)
);

NOR2_X4 _4934_ (
  .A1(\d_pipe[11][16] ),
  .A2(_0872_),
  .ZN(_0886_)
);

NAND2_X2 _4935_ (
  .A1(_0886_),
  .A2(_0880_),
  .ZN(_0887_)
);

NOR2_X4 _4936_ (
  .A1(_0887_),
  .A2(_0865_),
  .ZN(_0888_)
);

INV_X1 _4937_ (
  .A(\d_pipe[11][20] ),
  .ZN(_0889_)
);

XNOR2_X1 _4938_ (
  .A(_0888_),
  .B(_0889_),
  .ZN(_0890_)
);

OAI21_X1 _4939_ (
  .A(_0885_),
  .B1(_0890_),
  .B2(\s_pipe[11][24] ),
  .ZN(_4309_)
);

NAND4_X1 _4940_ (
  .A1(_0861_),
  .A2(_0869_),
  .A3(_0857_),
  .A4(_0858_),
  .ZN(_0891_)
);

NAND2_X1 _4941_ (
  .A1(_0873_),
  .A2(_0877_),
  .ZN(_0892_)
);

INV_X1 _4942_ (
  .A(\d_pipe[11][19] ),
  .ZN(_0893_)
);

NAND2_X1 _4943_ (
  .A1(_0893_),
  .A2(_0889_),
  .ZN(_0894_)
);

NOR3_X2 _4944_ (
  .A1(_0891_),
  .A2(_0892_),
  .A3(_0894_),
  .ZN(_0895_)
);

NAND2_X1 _4945_ (
  .A1(_0895_),
  .A2(_4285_),
  .ZN(_0896_)
);

NAND2_X1 _4946_ (
  .A1(_0896_),
  .A2(\d_pipe[11][21] ),
  .ZN(_0897_)
);

INV_X1 _4947_ (
  .A(\d_pipe[11][21] ),
  .ZN(_0898_)
);

NAND3_X1 _4948_ (
  .A1(_0895_),
  .A2(_4285_),
  .A3(_0898_),
  .ZN(_0899_)
);

NAND3_X1 _4949_ (
  .A1(_0897_),
  .A2(_0899_),
  .A3(_0637_),
  .ZN(_0900_)
);

OAI21_X1 _4950_ (
  .A(_0900_),
  .B1(_0855_),
  .B2(_0018_),
  .ZN(_4312_)
);

INV_X1 _4951_ (
  .A(_0888_),
  .ZN(_0901_)
);

NOR2_X2 _4952_ (
  .A1(\d_pipe[11][20] ),
  .A2(\d_pipe[11][21] ),
  .ZN(_0902_)
);

INV_X1 _4953_ (
  .A(\d_pipe[11][22] ),
  .ZN(_0903_)
);

NAND2_X1 _4954_ (
  .A1(_0902_),
  .A2(_0903_),
  .ZN(_0904_)
);

OAI21_X1 _4955_ (
  .A(_0637_),
  .B1(_0901_),
  .B2(_0904_),
  .ZN(_0905_)
);

AOI21_X1 _4956_ (
  .A(_0903_),
  .B1(_0888_),
  .B2(_0902_),
  .ZN(_0906_)
);

OAI22_X1 _4957_ (
  .A1(_0905_),
  .A2(_0906_),
  .B1(_0019_),
  .B2(_0855_),
  .ZN(_4315_)
);

NAND4_X1 _4958_ (
  .A1(_0898_),
  .A2(_0903_),
  .A3(_0893_),
  .A4(_0889_),
  .ZN(_0907_)
);

NOR2_X2 _4959_ (
  .A1(_0882_),
  .A2(_0907_),
  .ZN(_0908_)
);

INV_X1 _4960_ (
  .A(_0908_),
  .ZN(_0909_)
);

OAI21_X1 _4961_ (
  .A(\d_pipe[11][23] ),
  .B1(_0909_),
  .B2(_0859_),
  .ZN(_0910_)
);

INV_X1 _4962_ (
  .A(\d_pipe[11][23] ),
  .ZN(_0911_)
);

NAND3_X1 _4963_ (
  .A1(_0908_),
  .A2(_0911_),
  .A3(_0860_),
  .ZN(_0912_)
);

NAND3_X1 _4964_ (
  .A1(_0910_),
  .A2(_0637_),
  .A3(_0912_),
  .ZN(_0913_)
);

OAI21_X1 _4965_ (
  .A(_0913_),
  .B1(_0855_),
  .B2(_0020_),
  .ZN(_4318_)
);

XNOR2_X1 _4966_ (
  .A(_4323_),
  .B(\d_pipe[10][14] ),
  .ZN(_0914_)
);

BUF_X1 _4967_ (
  .A(_0638_),
  .Z(_0915_)
);

NAND2_X1 _4968_ (
  .A1(_0914_),
  .A2(_0915_),
  .ZN(_0916_)
);

OAI21_X1 _4969_ (
  .A(_0916_),
  .B1(_0915_),
  .B2(_0021_),
  .ZN(_4327_)
);

INV_X2 _4970_ (
  .A(\d_pipe[10][14] ),
  .ZN(_0917_)
);

INV_X1 _4971_ (
  .A(\d_pipe[10][13] ),
  .ZN(_0918_)
);

NAND3_X1 _4972_ (
  .A1(_0917_),
  .A2(_0918_),
  .A3(_4321_),
  .ZN(_0919_)
);

INV_X1 _4973_ (
  .A(_0919_),
  .ZN(_0920_)
);

INV_X4 _4974_ (
  .A(\d_pipe[10][15] ),
  .ZN(_0921_)
);

OAI21_X1 _4975_ (
  .A(_0639_),
  .B1(_0920_),
  .B2(_0921_),
  .ZN(_0922_)
);

NAND2_X1 _4976_ (
  .A1(_0920_),
  .A2(_0921_),
  .ZN(_0923_)
);

INV_X1 _4977_ (
  .A(_0923_),
  .ZN(_0924_)
);

OAI22_X1 _4978_ (
  .A1(_0922_),
  .A2(_0924_),
  .B1(_0022_),
  .B2(_0915_),
  .ZN(_4330_)
);

NAND3_X2 _4979_ (
  .A1(_0917_),
  .A2(_0921_),
  .A3(_4323_),
  .ZN(_0925_)
);

BUF_X4 _4980_ (
  .A(\d_pipe[10][16] ),
  .Z(_0926_)
);

OR2_X1 _4981_ (
  .A1(_0925_),
  .A2(_0926_),
  .ZN(_0927_)
);

NAND2_X1 _4982_ (
  .A1(_0925_),
  .A2(_0926_),
  .ZN(_0928_)
);

NAND3_X1 _4983_ (
  .A1(_0927_),
  .A2(_0639_),
  .A3(_0928_),
  .ZN(_0929_)
);

OAI21_X1 _4984_ (
  .A(_0929_),
  .B1(_0915_),
  .B2(_0023_),
  .ZN(_4333_)
);

INV_X2 _4985_ (
  .A(_0926_),
  .ZN(_0930_)
);

BUF_X4 _4986_ (
  .A(\d_pipe[10][17] ),
  .Z(_0931_)
);

INV_X2 _4987_ (
  .A(_0931_),
  .ZN(_0932_)
);

NAND3_X1 _4988_ (
  .A1(_0924_),
  .A2(_0930_),
  .A3(_0932_),
  .ZN(_0933_)
);

OAI21_X1 _4989_ (
  .A(_0931_),
  .B1(_0923_),
  .B2(_0926_),
  .ZN(_0934_)
);

NAND3_X1 _4990_ (
  .A1(_0933_),
  .A2(_0934_),
  .A3(_0639_),
  .ZN(_0935_)
);

OAI21_X1 _4991_ (
  .A(_0935_),
  .B1(_0915_),
  .B2(_0024_),
  .ZN(_4336_)
);

NOR2_X1 _4992_ (
  .A1(_0927_),
  .A2(_0931_),
  .ZN(_0936_)
);

INV_X1 _4993_ (
  .A(\d_pipe[10][18] ),
  .ZN(_0937_)
);

OAI21_X1 _4994_ (
  .A(_0639_),
  .B1(_0936_),
  .B2(_0937_),
  .ZN(_0938_)
);

NOR3_X1 _4995_ (
  .A1(_0927_),
  .A2(_0931_),
  .A3(\d_pipe[10][18] ),
  .ZN(_0939_)
);

OAI22_X1 _4996_ (
  .A1(_0938_),
  .A2(_0939_),
  .B1(_0025_),
  .B2(_0915_),
  .ZN(_4339_)
);

OR2_X1 _4997_ (
  .A1(_0639_),
  .A2(_0026_),
  .ZN(_0940_)
);

NAND4_X2 _4998_ (
  .A1(_0932_),
  .A2(_0937_),
  .A3(_0921_),
  .A4(_0930_),
  .ZN(_0941_)
);

NOR2_X1 _4999_ (
  .A1(_0941_),
  .A2(_0919_),
  .ZN(_0942_)
);

INV_X1 _5000_ (
  .A(\d_pipe[10][19] ),
  .ZN(_0943_)
);

XNOR2_X1 _5001_ (
  .A(_0942_),
  .B(_0943_),
  .ZN(_0944_)
);

OAI21_X1 _5002_ (
  .A(_0940_),
  .B1(_0944_),
  .B2(\s_pipe[10][24] ),
  .ZN(_4342_)
);

OR2_X1 _5003_ (
  .A1(_0639_),
  .A2(_0027_),
  .ZN(_0945_)
);

NOR2_X4 _5004_ (
  .A1(_0926_),
  .A2(_0931_),
  .ZN(_0946_)
);

NOR2_X1 _5005_ (
  .A1(\d_pipe[10][18] ),
  .A2(\d_pipe[10][19] ),
  .ZN(_0947_)
);

NAND2_X2 _5006_ (
  .A1(_0946_),
  .A2(_0947_),
  .ZN(_0948_)
);

NOR2_X4 _5007_ (
  .A1(_0948_),
  .A2(_0925_),
  .ZN(_0949_)
);

INV_X1 _5008_ (
  .A(\d_pipe[10][20] ),
  .ZN(_0950_)
);

XNOR2_X1 _5009_ (
  .A(_0949_),
  .B(_0950_),
  .ZN(_0951_)
);

OAI21_X1 _5010_ (
  .A(_0945_),
  .B1(_0951_),
  .B2(\s_pipe[10][24] ),
  .ZN(_4345_)
);

NAND4_X1 _5011_ (
  .A1(_0921_),
  .A2(_0930_),
  .A3(_0917_),
  .A4(_0918_),
  .ZN(_0952_)
);

NAND2_X1 _5012_ (
  .A1(_0932_),
  .A2(_0937_),
  .ZN(_0953_)
);

NAND2_X1 _5013_ (
  .A1(_0943_),
  .A2(_0950_),
  .ZN(_0954_)
);

NOR3_X2 _5014_ (
  .A1(_0952_),
  .A2(_0953_),
  .A3(_0954_),
  .ZN(_0955_)
);

NAND2_X1 _5015_ (
  .A1(_0955_),
  .A2(_4321_),
  .ZN(_0956_)
);

NAND2_X1 _5016_ (
  .A1(_0956_),
  .A2(\d_pipe[10][21] ),
  .ZN(_0957_)
);

INV_X1 _5017_ (
  .A(\d_pipe[10][21] ),
  .ZN(_0958_)
);

NAND3_X1 _5018_ (
  .A1(_0955_),
  .A2(_4321_),
  .A3(_0958_),
  .ZN(_0959_)
);

NAND3_X1 _5019_ (
  .A1(_0957_),
  .A2(_0959_),
  .A3(_0639_),
  .ZN(_0960_)
);

OAI21_X1 _5020_ (
  .A(_0960_),
  .B1(_0915_),
  .B2(_0028_),
  .ZN(_4348_)
);

INV_X1 _5021_ (
  .A(_0949_),
  .ZN(_0961_)
);

NOR2_X2 _5022_ (
  .A1(\d_pipe[10][20] ),
  .A2(\d_pipe[10][21] ),
  .ZN(_0962_)
);

INV_X1 _5023_ (
  .A(\d_pipe[10][22] ),
  .ZN(_0963_)
);

NAND2_X1 _5024_ (
  .A1(_0962_),
  .A2(_0963_),
  .ZN(_0964_)
);

OAI21_X1 _5025_ (
  .A(_0639_),
  .B1(_0961_),
  .B2(_0964_),
  .ZN(_0965_)
);

AOI21_X1 _5026_ (
  .A(_0963_),
  .B1(_0949_),
  .B2(_0962_),
  .ZN(_0966_)
);

OAI22_X1 _5027_ (
  .A1(_0965_),
  .A2(_0966_),
  .B1(_0029_),
  .B2(_0915_),
  .ZN(_4351_)
);

NAND4_X1 _5028_ (
  .A1(_0958_),
  .A2(_0963_),
  .A3(_0943_),
  .A4(_0950_),
  .ZN(_0967_)
);

NOR2_X1 _5029_ (
  .A1(_0941_),
  .A2(_0967_),
  .ZN(_0968_)
);

INV_X1 _5030_ (
  .A(_0968_),
  .ZN(_0969_)
);

OAI21_X1 _5031_ (
  .A(\d_pipe[10][23] ),
  .B1(_0969_),
  .B2(_0919_),
  .ZN(_0970_)
);

INV_X1 _5032_ (
  .A(\d_pipe[10][23] ),
  .ZN(_0971_)
);

NAND3_X1 _5033_ (
  .A1(_0968_),
  .A2(_0971_),
  .A3(_0920_),
  .ZN(_0972_)
);

NAND3_X1 _5034_ (
  .A1(_0970_),
  .A2(_0915_),
  .A3(_0972_),
  .ZN(_0973_)
);

OAI21_X1 _5035_ (
  .A(_0973_),
  .B1(_0915_),
  .B2(_0030_),
  .ZN(_4354_)
);

AOI21_X1 _5036_ (
  .A(_0641_),
  .B1(_0679_),
  .B2(_4359_),
  .ZN(_0974_)
);

OAI21_X1 _5037_ (
  .A(_0974_),
  .B1(_4359_),
  .B2(_0679_),
  .ZN(_0975_)
);

OAI21_X1 _5038_ (
  .A(_0975_),
  .B1(_0684_),
  .B2(_0031_),
  .ZN(_4363_)
);

INV_X1 _5039_ (
  .A(_3714_),
  .ZN(_0976_)
);

NAND3_X1 _5040_ (
  .A1(_0679_),
  .A2(_0976_),
  .A3(_4357_),
  .ZN(_0977_)
);

INV_X1 _5041_ (
  .A(_0977_),
  .ZN(_0978_)
);

OAI21_X1 _5042_ (
  .A(_0643_),
  .B1(_0978_),
  .B2(_0680_),
  .ZN(_0979_)
);

NAND2_X1 _5043_ (
  .A1(_0978_),
  .A2(_0680_),
  .ZN(_0980_)
);

INV_X1 _5044_ (
  .A(_0980_),
  .ZN(_0981_)
);

OAI22_X1 _5045_ (
  .A1(_0979_),
  .A2(_0981_),
  .B1(_0032_),
  .B2(_0684_),
  .ZN(_4366_)
);

INV_X2 _5046_ (
  .A(_0682_),
  .ZN(_0982_)
);

BUF_X4 _5047_ (
  .A(_3718_),
  .Z(_0983_)
);

INV_X2 _5048_ (
  .A(_0983_),
  .ZN(_0984_)
);

NAND3_X1 _5049_ (
  .A1(_0981_),
  .A2(_0982_),
  .A3(_0984_),
  .ZN(_0985_)
);

OAI21_X1 _5050_ (
  .A(_0983_),
  .B1(_0980_),
  .B2(_0682_),
  .ZN(_0986_)
);

NAND3_X1 _5051_ (
  .A1(_0985_),
  .A2(_0986_),
  .A3(_0643_),
  .ZN(_0987_)
);

OAI21_X1 _5052_ (
  .A(_0987_),
  .B1(_0684_),
  .B2(_0034_),
  .ZN(_4372_)
);

NOR2_X1 _5053_ (
  .A1(_0683_),
  .A2(_0983_),
  .ZN(_0988_)
);

INV_X1 _5054_ (
  .A(_3719_),
  .ZN(_0989_)
);

OAI21_X1 _5055_ (
  .A(_0643_),
  .B1(_0988_),
  .B2(_0989_),
  .ZN(_0990_)
);

NOR3_X1 _5056_ (
  .A1(_0683_),
  .A2(_0983_),
  .A3(_3719_),
  .ZN(_0991_)
);

OAI22_X1 _5057_ (
  .A1(_0990_),
  .A2(_0991_),
  .B1(_0035_),
  .B2(_0684_),
  .ZN(_4375_)
);

OR2_X1 _5058_ (
  .A1(_0643_),
  .A2(_0036_),
  .ZN(_0992_)
);

NAND4_X2 _5059_ (
  .A1(_0984_),
  .A2(_0989_),
  .A3(_0680_),
  .A4(_0982_),
  .ZN(_0993_)
);

NOR2_X1 _5060_ (
  .A1(_0993_),
  .A2(_0977_),
  .ZN(_0994_)
);

INV_X1 _5061_ (
  .A(_3720_),
  .ZN(_0995_)
);

XNOR2_X1 _5062_ (
  .A(_0994_),
  .B(_0995_),
  .ZN(_0996_)
);

OAI21_X1 _5063_ (
  .A(_0992_),
  .B1(_0996_),
  .B2(_0641_),
  .ZN(_4378_)
);

OR2_X1 _5064_ (
  .A1(_0643_),
  .A2(_0037_),
  .ZN(_0997_)
);

NOR2_X4 _5065_ (
  .A1(_0682_),
  .A2(_0983_),
  .ZN(_0998_)
);

NOR2_X1 _5066_ (
  .A1(_3719_),
  .A2(_3720_),
  .ZN(_0999_)
);

NAND2_X2 _5067_ (
  .A1(_0998_),
  .A2(_0999_),
  .ZN(_1000_)
);

NOR2_X4 _5068_ (
  .A1(_1000_),
  .A2(_0681_),
  .ZN(_1001_)
);

INV_X1 _5069_ (
  .A(_3721_),
  .ZN(_1002_)
);

XNOR2_X1 _5070_ (
  .A(_1001_),
  .B(_1002_),
  .ZN(_1003_)
);

OAI21_X1 _5071_ (
  .A(_0997_),
  .B1(_1003_),
  .B2(_0641_),
  .ZN(_4381_)
);

NAND4_X1 _5072_ (
  .A1(_0680_),
  .A2(_0982_),
  .A3(_0679_),
  .A4(_0976_),
  .ZN(_1004_)
);

NAND2_X1 _5073_ (
  .A1(_0984_),
  .A2(_0989_),
  .ZN(_1005_)
);

NAND2_X1 _5074_ (
  .A1(_0995_),
  .A2(_1002_),
  .ZN(_1006_)
);

NOR3_X2 _5075_ (
  .A1(_1004_),
  .A2(_1005_),
  .A3(_1006_),
  .ZN(_1007_)
);

NAND2_X1 _5076_ (
  .A1(_1007_),
  .A2(_4357_),
  .ZN(_1008_)
);

NAND2_X1 _5077_ (
  .A1(_1008_),
  .A2(_3722_),
  .ZN(_1009_)
);

INV_X1 _5078_ (
  .A(_3722_),
  .ZN(_1010_)
);

NAND3_X1 _5079_ (
  .A1(_1007_),
  .A2(_4357_),
  .A3(_1010_),
  .ZN(_1011_)
);

NAND3_X1 _5080_ (
  .A1(_1009_),
  .A2(_1011_),
  .A3(_0643_),
  .ZN(_1012_)
);

OAI21_X1 _5081_ (
  .A(_1012_),
  .B1(_0684_),
  .B2(_0038_),
  .ZN(_4384_)
);

INV_X1 _5082_ (
  .A(_1001_),
  .ZN(_1013_)
);

NOR2_X2 _5083_ (
  .A1(_3721_),
  .A2(_3722_),
  .ZN(_1014_)
);

INV_X1 _5084_ (
  .A(_3712_),
  .ZN(_1015_)
);

NAND2_X1 _5085_ (
  .A1(_1014_),
  .A2(_1015_),
  .ZN(_1016_)
);

OAI21_X1 _5086_ (
  .A(_0643_),
  .B1(_1013_),
  .B2(_1016_),
  .ZN(_1017_)
);

AOI21_X1 _5087_ (
  .A(_1015_),
  .B1(_1001_),
  .B2(_1014_),
  .ZN(_1018_)
);

OAI22_X1 _5088_ (
  .A1(_1017_),
  .A2(_1018_),
  .B1(_0039_),
  .B2(_0684_),
  .ZN(_4387_)
);

NAND4_X1 _5089_ (
  .A1(_1010_),
  .A2(_1015_),
  .A3(_0995_),
  .A4(_1002_),
  .ZN(_1019_)
);

NOR2_X2 _5090_ (
  .A1(_0993_),
  .A2(_1019_),
  .ZN(_1020_)
);

INV_X1 _5091_ (
  .A(_1020_),
  .ZN(_1021_)
);

OAI21_X1 _5092_ (
  .A(_3713_),
  .B1(_1021_),
  .B2(_0977_),
  .ZN(_1022_)
);

INV_X1 _5093_ (
  .A(_3713_),
  .ZN(_1023_)
);

NAND3_X1 _5094_ (
  .A1(_1020_),
  .A2(_1023_),
  .A3(_0978_),
  .ZN(_1024_)
);

NAND3_X1 _5095_ (
  .A1(_1022_),
  .A2(_0684_),
  .A3(_1024_),
  .ZN(_1025_)
);

OAI21_X1 _5096_ (
  .A(_1025_),
  .B1(_0684_),
  .B2(_0040_),
  .ZN(_4390_)
);

XNOR2_X1 _5097_ (
  .A(_4395_),
  .B(\d_pipe[8][14] ),
  .ZN(_1026_)
);

BUF_X1 _5098_ (
  .A(_0645_),
  .Z(_1027_)
);

NAND2_X1 _5099_ (
  .A1(_1026_),
  .A2(_1027_),
  .ZN(_1028_)
);

OAI21_X1 _5100_ (
  .A(_1028_),
  .B1(_1027_),
  .B2(_0041_),
  .ZN(_4399_)
);

INV_X2 _5101_ (
  .A(\d_pipe[8][14] ),
  .ZN(_1029_)
);

INV_X1 _5102_ (
  .A(\d_pipe[8][13] ),
  .ZN(_1030_)
);

NAND3_X2 _5103_ (
  .A1(_1029_),
  .A2(_1030_),
  .A3(_4393_),
  .ZN(_1031_)
);

INV_X2 _5104_ (
  .A(_1031_),
  .ZN(_1032_)
);

INV_X4 _5105_ (
  .A(\d_pipe[8][15] ),
  .ZN(_1033_)
);

OAI21_X1 _5106_ (
  .A(_0647_),
  .B1(_1032_),
  .B2(_1033_),
  .ZN(_1034_)
);

NAND2_X1 _5107_ (
  .A1(_1032_),
  .A2(_1033_),
  .ZN(_1035_)
);

INV_X2 _5108_ (
  .A(_1035_),
  .ZN(_1036_)
);

OAI22_X1 _5109_ (
  .A1(_1034_),
  .A2(_1036_),
  .B1(_0042_),
  .B2(_1027_),
  .ZN(_4402_)
);

NAND3_X2 _5110_ (
  .A1(_1029_),
  .A2(_1033_),
  .A3(_4395_),
  .ZN(_1037_)
);

BUF_X2 _5111_ (
  .A(\d_pipe[8][16] ),
  .Z(_1038_)
);

OR2_X1 _5112_ (
  .A1(_1037_),
  .A2(_1038_),
  .ZN(_1039_)
);

NAND2_X1 _5113_ (
  .A1(_1037_),
  .A2(_1038_),
  .ZN(_1040_)
);

NAND3_X1 _5114_ (
  .A1(_1039_),
  .A2(_0647_),
  .A3(_1040_),
  .ZN(_1041_)
);

OAI21_X1 _5115_ (
  .A(_1041_),
  .B1(_1027_),
  .B2(_0043_),
  .ZN(_4405_)
);

INV_X4 _5116_ (
  .A(_1038_),
  .ZN(_1042_)
);

NAND2_X1 _5117_ (
  .A1(_1036_),
  .A2(_1042_),
  .ZN(_1043_)
);

INV_X1 _5118_ (
  .A(_1043_),
  .ZN(_1044_)
);

BUF_X4 _5119_ (
  .A(\d_pipe[8][17] ),
  .Z(_1045_)
);

INV_X2 _5120_ (
  .A(_1045_),
  .ZN(_1046_)
);

OAI21_X1 _5121_ (
  .A(_0647_),
  .B1(_1044_),
  .B2(_1046_),
  .ZN(_1047_)
);

NOR2_X2 _5122_ (
  .A1(_1043_),
  .A2(_1045_),
  .ZN(_1048_)
);

OAI22_X1 _5123_ (
  .A1(_1047_),
  .A2(_1048_),
  .B1(_0044_),
  .B2(_1027_),
  .ZN(_4408_)
);

NOR2_X1 _5124_ (
  .A1(_1039_),
  .A2(_1045_),
  .ZN(_1049_)
);

INV_X1 _5125_ (
  .A(\d_pipe[8][18] ),
  .ZN(_1050_)
);

OAI21_X1 _5126_ (
  .A(_0647_),
  .B1(_1049_),
  .B2(_1050_),
  .ZN(_1051_)
);

NOR3_X1 _5127_ (
  .A1(_1039_),
  .A2(_1045_),
  .A3(\d_pipe[8][18] ),
  .ZN(_1052_)
);

OAI22_X1 _5128_ (
  .A1(_1051_),
  .A2(_1052_),
  .B1(_0045_),
  .B2(_1027_),
  .ZN(_4411_)
);

NOR2_X2 _5129_ (
  .A1(\d_pipe[8][18] ),
  .A2(\d_pipe[8][19] ),
  .ZN(_1053_)
);

NAND2_X1 _5130_ (
  .A1(_1048_),
  .A2(_1053_),
  .ZN(_1054_)
);

NAND4_X2 _5131_ (
  .A1(_1046_),
  .A2(_1050_),
  .A3(_1033_),
  .A4(_1042_),
  .ZN(_1055_)
);

OAI21_X1 _5132_ (
  .A(\d_pipe[8][19] ),
  .B1(_1055_),
  .B2(_1031_),
  .ZN(_1056_)
);

NAND3_X1 _5133_ (
  .A1(_1054_),
  .A2(_0647_),
  .A3(_1056_),
  .ZN(_1057_)
);

OAI21_X1 _5134_ (
  .A(_1057_),
  .B1(_1027_),
  .B2(_0046_),
  .ZN(_4414_)
);

OR2_X1 _5135_ (
  .A1(_0647_),
  .A2(_0047_),
  .ZN(_1058_)
);

NOR2_X4 _5136_ (
  .A1(_1038_),
  .A2(_1045_),
  .ZN(_1059_)
);

NAND2_X2 _5137_ (
  .A1(_1059_),
  .A2(_1053_),
  .ZN(_1060_)
);

NOR2_X4 _5138_ (
  .A1(_1060_),
  .A2(_1037_),
  .ZN(_1061_)
);

INV_X1 _5139_ (
  .A(\d_pipe[8][20] ),
  .ZN(_1062_)
);

XNOR2_X1 _5140_ (
  .A(_1061_),
  .B(_1062_),
  .ZN(_1063_)
);

OAI21_X1 _5141_ (
  .A(_1058_),
  .B1(_1063_),
  .B2(\s_pipe[8][24] ),
  .ZN(_4417_)
);

NAND4_X1 _5142_ (
  .A1(_1033_),
  .A2(_1042_),
  .A3(_1029_),
  .A4(_1030_),
  .ZN(_1064_)
);

NAND2_X1 _5143_ (
  .A1(_1046_),
  .A2(_1050_),
  .ZN(_1065_)
);

INV_X1 _5144_ (
  .A(\d_pipe[8][19] ),
  .ZN(_1066_)
);

NAND2_X1 _5145_ (
  .A1(_1066_),
  .A2(_1062_),
  .ZN(_1067_)
);

NOR3_X2 _5146_ (
  .A1(_1064_),
  .A2(_1065_),
  .A3(_1067_),
  .ZN(_1068_)
);

NAND2_X1 _5147_ (
  .A1(_1068_),
  .A2(_4393_),
  .ZN(_1069_)
);

NAND2_X1 _5148_ (
  .A1(_1069_),
  .A2(\d_pipe[8][21] ),
  .ZN(_1070_)
);

INV_X1 _5149_ (
  .A(\d_pipe[8][21] ),
  .ZN(_1071_)
);

NAND3_X1 _5150_ (
  .A1(_1068_),
  .A2(_4393_),
  .A3(_1071_),
  .ZN(_1072_)
);

NAND3_X1 _5151_ (
  .A1(_1070_),
  .A2(_1072_),
  .A3(_0647_),
  .ZN(_1073_)
);

OAI21_X1 _5152_ (
  .A(_1073_),
  .B1(_1027_),
  .B2(_0048_),
  .ZN(_4420_)
);

INV_X1 _5153_ (
  .A(_1061_),
  .ZN(_1074_)
);

NOR2_X2 _5154_ (
  .A1(\d_pipe[8][20] ),
  .A2(\d_pipe[8][21] ),
  .ZN(_1075_)
);

INV_X1 _5155_ (
  .A(\d_pipe[8][22] ),
  .ZN(_1076_)
);

NAND2_X1 _5156_ (
  .A1(_1075_),
  .A2(_1076_),
  .ZN(_1077_)
);

OAI21_X1 _5157_ (
  .A(_0647_),
  .B1(_1074_),
  .B2(_1077_),
  .ZN(_1078_)
);

AOI21_X1 _5158_ (
  .A(_1076_),
  .B1(_1061_),
  .B2(_1075_),
  .ZN(_1079_)
);

OAI22_X1 _5159_ (
  .A1(_1078_),
  .A2(_1079_),
  .B1(_0049_),
  .B2(_1027_),
  .ZN(_4423_)
);

NAND4_X1 _5160_ (
  .A1(_1071_),
  .A2(_1076_),
  .A3(_1066_),
  .A4(_1062_),
  .ZN(_1080_)
);

NOR2_X2 _5161_ (
  .A1(_1055_),
  .A2(_1080_),
  .ZN(_1081_)
);

INV_X1 _5162_ (
  .A(_1081_),
  .ZN(_1082_)
);

OAI21_X1 _5163_ (
  .A(\d_pipe[8][23] ),
  .B1(_1082_),
  .B2(_1031_),
  .ZN(_1083_)
);

INV_X1 _5164_ (
  .A(\d_pipe[8][23] ),
  .ZN(_1084_)
);

NAND3_X1 _5165_ (
  .A1(_1081_),
  .A2(_1084_),
  .A3(_1032_),
  .ZN(_1085_)
);

NAND3_X1 _5166_ (
  .A1(_1083_),
  .A2(_0647_),
  .A3(_1085_),
  .ZN(_1086_)
);

OAI21_X1 _5167_ (
  .A(_1086_),
  .B1(_1027_),
  .B2(_0050_),
  .ZN(_4426_)
);

XNOR2_X1 _5168_ (
  .A(_4431_),
  .B(\d_pipe[7][14] ),
  .ZN(_1087_)
);

BUF_X1 _5169_ (
  .A(_0648_),
  .Z(_1088_)
);

NAND2_X1 _5170_ (
  .A1(_1087_),
  .A2(_1088_),
  .ZN(_1089_)
);

OAI21_X1 _5171_ (
  .A(_1089_),
  .B1(_1088_),
  .B2(_0051_),
  .ZN(_4435_)
);

INV_X2 _5172_ (
  .A(\d_pipe[7][14] ),
  .ZN(_1090_)
);

INV_X2 _5173_ (
  .A(\d_pipe[7][13] ),
  .ZN(_1091_)
);

NAND3_X2 _5174_ (
  .A1(_1090_),
  .A2(_1091_),
  .A3(_4429_),
  .ZN(_1092_)
);

INV_X2 _5175_ (
  .A(_1092_),
  .ZN(_1093_)
);

INV_X4 _5176_ (
  .A(\d_pipe[7][15] ),
  .ZN(_1094_)
);

OAI21_X1 _5177_ (
  .A(_0650_),
  .B1(_1093_),
  .B2(_1094_),
  .ZN(_1095_)
);

NAND2_X1 _5178_ (
  .A1(_1093_),
  .A2(_1094_),
  .ZN(_1096_)
);

INV_X1 _5179_ (
  .A(_1096_),
  .ZN(_1097_)
);

OAI22_X1 _5180_ (
  .A1(_1095_),
  .A2(_1097_),
  .B1(_0052_),
  .B2(_1088_),
  .ZN(_4438_)
);

NAND3_X2 _5181_ (
  .A1(_1090_),
  .A2(_1094_),
  .A3(_4431_),
  .ZN(_1098_)
);

BUF_X4 _5182_ (
  .A(\d_pipe[7][16] ),
  .Z(_1099_)
);

OR2_X1 _5183_ (
  .A1(_1098_),
  .A2(_1099_),
  .ZN(_1100_)
);

NAND2_X1 _5184_ (
  .A1(_1098_),
  .A2(_1099_),
  .ZN(_1101_)
);

NAND3_X1 _5185_ (
  .A1(_1100_),
  .A2(_0650_),
  .A3(_1101_),
  .ZN(_1102_)
);

OAI21_X1 _5186_ (
  .A(_1102_),
  .B1(_1088_),
  .B2(_0053_),
  .ZN(_4441_)
);

INV_X2 _5187_ (
  .A(_1099_),
  .ZN(_1103_)
);

NAND2_X1 _5188_ (
  .A1(_1097_),
  .A2(_1103_),
  .ZN(_1104_)
);

INV_X1 _5189_ (
  .A(_1104_),
  .ZN(_1105_)
);

BUF_X4 _5190_ (
  .A(\d_pipe[7][17] ),
  .Z(_1106_)
);

INV_X2 _5191_ (
  .A(_1106_),
  .ZN(_1107_)
);

OAI21_X1 _5192_ (
  .A(_0650_),
  .B1(_1105_),
  .B2(_1107_),
  .ZN(_1108_)
);

NOR2_X2 _5193_ (
  .A1(_1104_),
  .A2(_1106_),
  .ZN(_1109_)
);

OAI22_X1 _5194_ (
  .A1(_1108_),
  .A2(_1109_),
  .B1(_0054_),
  .B2(_1088_),
  .ZN(_4444_)
);

NOR2_X1 _5195_ (
  .A1(_1100_),
  .A2(_1106_),
  .ZN(_1110_)
);

INV_X1 _5196_ (
  .A(\d_pipe[7][18] ),
  .ZN(_1111_)
);

OAI21_X1 _5197_ (
  .A(_0650_),
  .B1(_1110_),
  .B2(_1111_),
  .ZN(_1112_)
);

NOR3_X1 _5198_ (
  .A1(_1100_),
  .A2(_1106_),
  .A3(\d_pipe[7][18] ),
  .ZN(_1113_)
);

OAI22_X1 _5199_ (
  .A1(_1112_),
  .A2(_1113_),
  .B1(_0055_),
  .B2(_1088_),
  .ZN(_4447_)
);

NOR2_X2 _5200_ (
  .A1(\d_pipe[7][18] ),
  .A2(\d_pipe[7][19] ),
  .ZN(_1114_)
);

NAND2_X1 _5201_ (
  .A1(_1109_),
  .A2(_1114_),
  .ZN(_1115_)
);

NAND4_X2 _5202_ (
  .A1(_1107_),
  .A2(_1111_),
  .A3(_1094_),
  .A4(_1103_),
  .ZN(_1116_)
);

OAI21_X1 _5203_ (
  .A(\d_pipe[7][19] ),
  .B1(_1116_),
  .B2(_1092_),
  .ZN(_1117_)
);

NAND3_X1 _5204_ (
  .A1(_1115_),
  .A2(_0650_),
  .A3(_1117_),
  .ZN(_1118_)
);

OAI21_X1 _5205_ (
  .A(_1118_),
  .B1(_1088_),
  .B2(_0056_),
  .ZN(_4450_)
);

OR2_X1 _5206_ (
  .A1(_0650_),
  .A2(_0057_),
  .ZN(_1119_)
);

NOR2_X4 _5207_ (
  .A1(_1099_),
  .A2(_1106_),
  .ZN(_1120_)
);

NAND2_X2 _5208_ (
  .A1(_1120_),
  .A2(_1114_),
  .ZN(_1121_)
);

NOR2_X4 _5209_ (
  .A1(_1121_),
  .A2(_1098_),
  .ZN(_1122_)
);

INV_X1 _5210_ (
  .A(\d_pipe[7][20] ),
  .ZN(_1123_)
);

XNOR2_X1 _5211_ (
  .A(_1122_),
  .B(_1123_),
  .ZN(_1124_)
);

OAI21_X1 _5212_ (
  .A(_1119_),
  .B1(_1124_),
  .B2(\s_pipe[7][24] ),
  .ZN(_4453_)
);

NAND4_X1 _5213_ (
  .A1(_1094_),
  .A2(_1103_),
  .A3(_1090_),
  .A4(_1091_),
  .ZN(_1125_)
);

NAND2_X1 _5214_ (
  .A1(_1107_),
  .A2(_1111_),
  .ZN(_1126_)
);

INV_X1 _5215_ (
  .A(\d_pipe[7][19] ),
  .ZN(_1127_)
);

NAND2_X1 _5216_ (
  .A1(_1127_),
  .A2(_1123_),
  .ZN(_1128_)
);

NOR3_X2 _5217_ (
  .A1(_1125_),
  .A2(_1126_),
  .A3(_1128_),
  .ZN(_1129_)
);

NAND2_X1 _5218_ (
  .A1(_1129_),
  .A2(_4429_),
  .ZN(_1130_)
);

NAND2_X1 _5219_ (
  .A1(_1130_),
  .A2(\d_pipe[7][21] ),
  .ZN(_1131_)
);

INV_X1 _5220_ (
  .A(\d_pipe[7][21] ),
  .ZN(_1132_)
);

NAND3_X1 _5221_ (
  .A1(_1129_),
  .A2(_4429_),
  .A3(_1132_),
  .ZN(_1133_)
);

NAND3_X1 _5222_ (
  .A1(_1131_),
  .A2(_1133_),
  .A3(_0650_),
  .ZN(_1134_)
);

OAI21_X1 _5223_ (
  .A(_1134_),
  .B1(_1088_),
  .B2(_0058_),
  .ZN(_4456_)
);

INV_X1 _5224_ (
  .A(_1122_),
  .ZN(_1135_)
);

NOR2_X2 _5225_ (
  .A1(\d_pipe[7][20] ),
  .A2(\d_pipe[7][21] ),
  .ZN(_1136_)
);

INV_X1 _5226_ (
  .A(\d_pipe[7][22] ),
  .ZN(_1137_)
);

NAND2_X1 _5227_ (
  .A1(_1136_),
  .A2(_1137_),
  .ZN(_1138_)
);

OAI21_X1 _5228_ (
  .A(_0650_),
  .B1(_1135_),
  .B2(_1138_),
  .ZN(_1139_)
);

AOI21_X1 _5229_ (
  .A(_1137_),
  .B1(_1122_),
  .B2(_1136_),
  .ZN(_1140_)
);

OAI22_X1 _5230_ (
  .A1(_1139_),
  .A2(_1140_),
  .B1(_0059_),
  .B2(_1088_),
  .ZN(_4459_)
);

NAND4_X1 _5231_ (
  .A1(_1132_),
  .A2(_1137_),
  .A3(_1127_),
  .A4(_1123_),
  .ZN(_1141_)
);

NOR2_X1 _5232_ (
  .A1(_1116_),
  .A2(_1141_),
  .ZN(_1142_)
);

INV_X1 _5233_ (
  .A(_1142_),
  .ZN(_1143_)
);

OAI21_X1 _5234_ (
  .A(\d_pipe[7][23] ),
  .B1(_1143_),
  .B2(_1092_),
  .ZN(_1144_)
);

INV_X1 _5235_ (
  .A(\d_pipe[7][23] ),
  .ZN(_1145_)
);

NAND3_X1 _5236_ (
  .A1(_1142_),
  .A2(_1145_),
  .A3(_1093_),
  .ZN(_1146_)
);

NAND3_X1 _5237_ (
  .A1(_1144_),
  .A2(_0650_),
  .A3(_1146_),
  .ZN(_1147_)
);

OAI21_X1 _5238_ (
  .A(_1147_),
  .B1(_1088_),
  .B2(_0060_),
  .ZN(_4462_)
);

XNOR2_X1 _5239_ (
  .A(_4467_),
  .B(\d_pipe[6][14] ),
  .ZN(_1148_)
);

BUF_X1 _5240_ (
  .A(_0651_),
  .Z(_1149_)
);

NAND2_X1 _5241_ (
  .A1(_1148_),
  .A2(_1149_),
  .ZN(_1150_)
);

OAI21_X1 _5242_ (
  .A(_1150_),
  .B1(_1149_),
  .B2(_0061_),
  .ZN(_4471_)
);

INV_X2 _5243_ (
  .A(\d_pipe[6][14] ),
  .ZN(_1151_)
);

INV_X1 _5244_ (
  .A(\d_pipe[6][13] ),
  .ZN(_1152_)
);

NAND3_X1 _5245_ (
  .A1(_1151_),
  .A2(_1152_),
  .A3(_4465_),
  .ZN(_1153_)
);

INV_X1 _5246_ (
  .A(_1153_),
  .ZN(_1154_)
);

INV_X2 _5247_ (
  .A(\d_pipe[6][15] ),
  .ZN(_1155_)
);

OAI21_X1 _5248_ (
  .A(_0652_),
  .B1(_1154_),
  .B2(_1155_),
  .ZN(_1156_)
);

NAND2_X1 _5249_ (
  .A1(_1154_),
  .A2(_1155_),
  .ZN(_1157_)
);

INV_X1 _5250_ (
  .A(_1157_),
  .ZN(_1158_)
);

OAI22_X1 _5251_ (
  .A1(_1156_),
  .A2(_1158_),
  .B1(_0062_),
  .B2(_1149_),
  .ZN(_4474_)
);

NAND3_X2 _5252_ (
  .A1(_1151_),
  .A2(_1155_),
  .A3(_4467_),
  .ZN(_1159_)
);

BUF_X4 _5253_ (
  .A(\d_pipe[6][16] ),
  .Z(_1160_)
);

OR2_X1 _5254_ (
  .A1(_1159_),
  .A2(_1160_),
  .ZN(_1161_)
);

NAND2_X1 _5255_ (
  .A1(_1159_),
  .A2(_1160_),
  .ZN(_1162_)
);

NAND3_X1 _5256_ (
  .A1(_1161_),
  .A2(_0652_),
  .A3(_1162_),
  .ZN(_1163_)
);

OAI21_X1 _5257_ (
  .A(_1163_),
  .B1(_1149_),
  .B2(_0063_),
  .ZN(_4477_)
);

INV_X4 _5258_ (
  .A(_1160_),
  .ZN(_1164_)
);

BUF_X4 _5259_ (
  .A(\d_pipe[6][17] ),
  .Z(_1165_)
);

INV_X2 _5260_ (
  .A(_1165_),
  .ZN(_1166_)
);

NAND3_X1 _5261_ (
  .A1(_1158_),
  .A2(_1164_),
  .A3(_1166_),
  .ZN(_1167_)
);

OAI21_X1 _5262_ (
  .A(_1165_),
  .B1(_1157_),
  .B2(_1160_),
  .ZN(_1168_)
);

NAND3_X1 _5263_ (
  .A1(_1167_),
  .A2(_1168_),
  .A3(_0652_),
  .ZN(_1169_)
);

OAI21_X1 _5264_ (
  .A(_1169_),
  .B1(_1149_),
  .B2(_0064_),
  .ZN(_4480_)
);

NOR2_X1 _5265_ (
  .A1(_1161_),
  .A2(_1165_),
  .ZN(_1170_)
);

INV_X1 _5266_ (
  .A(\d_pipe[6][18] ),
  .ZN(_1171_)
);

OAI21_X1 _5267_ (
  .A(_0652_),
  .B1(_1170_),
  .B2(_1171_),
  .ZN(_1172_)
);

NOR3_X1 _5268_ (
  .A1(_1161_),
  .A2(_1165_),
  .A3(\d_pipe[6][18] ),
  .ZN(_1173_)
);

OAI22_X1 _5269_ (
  .A1(_1172_),
  .A2(_1173_),
  .B1(_0065_),
  .B2(_1149_),
  .ZN(_4483_)
);

OR2_X1 _5270_ (
  .A1(_0652_),
  .A2(_0066_),
  .ZN(_1174_)
);

NAND4_X1 _5271_ (
  .A1(_1166_),
  .A2(_1171_),
  .A3(_1155_),
  .A4(_1164_),
  .ZN(_1175_)
);

NOR2_X1 _5272_ (
  .A1(_1175_),
  .A2(_1153_),
  .ZN(_1176_)
);

INV_X1 _5273_ (
  .A(\d_pipe[6][19] ),
  .ZN(_1177_)
);

XNOR2_X1 _5274_ (
  .A(_1176_),
  .B(_1177_),
  .ZN(_1178_)
);

OAI21_X1 _5275_ (
  .A(_1174_),
  .B1(_1178_),
  .B2(\s_pipe[6][24] ),
  .ZN(_4486_)
);

OR2_X1 _5276_ (
  .A1(_0652_),
  .A2(_0067_),
  .ZN(_1179_)
);

NOR2_X2 _5277_ (
  .A1(_1160_),
  .A2(_1165_),
  .ZN(_1180_)
);

NOR2_X1 _5278_ (
  .A1(\d_pipe[6][18] ),
  .A2(\d_pipe[6][19] ),
  .ZN(_1181_)
);

NAND2_X2 _5279_ (
  .A1(_1180_),
  .A2(_1181_),
  .ZN(_1182_)
);

NOR2_X4 _5280_ (
  .A1(_1182_),
  .A2(_1159_),
  .ZN(_1183_)
);

INV_X1 _5281_ (
  .A(\d_pipe[6][20] ),
  .ZN(_1184_)
);

XNOR2_X1 _5282_ (
  .A(_1183_),
  .B(_1184_),
  .ZN(_1185_)
);

OAI21_X1 _5283_ (
  .A(_1179_),
  .B1(_1185_),
  .B2(\s_pipe[6][24] ),
  .ZN(_4489_)
);

NAND4_X1 _5284_ (
  .A1(_1155_),
  .A2(_1164_),
  .A3(_1151_),
  .A4(_1152_),
  .ZN(_1186_)
);

NAND2_X1 _5285_ (
  .A1(_1166_),
  .A2(_1171_),
  .ZN(_1187_)
);

NAND2_X1 _5286_ (
  .A1(_1177_),
  .A2(_1184_),
  .ZN(_1188_)
);

NOR3_X2 _5287_ (
  .A1(_1186_),
  .A2(_1187_),
  .A3(_1188_),
  .ZN(_1189_)
);

NAND2_X1 _5288_ (
  .A1(_1189_),
  .A2(_4465_),
  .ZN(_1190_)
);

NAND2_X1 _5289_ (
  .A1(_1190_),
  .A2(\d_pipe[6][21] ),
  .ZN(_1191_)
);

INV_X1 _5290_ (
  .A(\d_pipe[6][21] ),
  .ZN(_1192_)
);

NAND3_X1 _5291_ (
  .A1(_1189_),
  .A2(_4465_),
  .A3(_1192_),
  .ZN(_1193_)
);

NAND3_X1 _5292_ (
  .A1(_1191_),
  .A2(_1193_),
  .A3(_0652_),
  .ZN(_1194_)
);

OAI21_X1 _5293_ (
  .A(_1194_),
  .B1(_1149_),
  .B2(_0068_),
  .ZN(_4492_)
);

INV_X1 _5294_ (
  .A(_1183_),
  .ZN(_1195_)
);

NOR2_X2 _5295_ (
  .A1(\d_pipe[6][20] ),
  .A2(\d_pipe[6][21] ),
  .ZN(_1196_)
);

INV_X1 _5296_ (
  .A(\d_pipe[6][22] ),
  .ZN(_1197_)
);

NAND2_X1 _5297_ (
  .A1(_1196_),
  .A2(_1197_),
  .ZN(_1198_)
);

OAI21_X1 _5298_ (
  .A(_0652_),
  .B1(_1195_),
  .B2(_1198_),
  .ZN(_1199_)
);

AOI21_X1 _5299_ (
  .A(_1197_),
  .B1(_1183_),
  .B2(_1196_),
  .ZN(_1200_)
);

OAI22_X1 _5300_ (
  .A1(_1199_),
  .A2(_1200_),
  .B1(_0069_),
  .B2(_1149_),
  .ZN(_4495_)
);

NAND4_X1 _5301_ (
  .A1(_1192_),
  .A2(_1197_),
  .A3(_1177_),
  .A4(_1184_),
  .ZN(_1201_)
);

NOR2_X1 _5302_ (
  .A1(_1175_),
  .A2(_1201_),
  .ZN(_1202_)
);

INV_X1 _5303_ (
  .A(_1202_),
  .ZN(_1203_)
);

OAI21_X1 _5304_ (
  .A(\d_pipe[6][23] ),
  .B1(_1203_),
  .B2(_1153_),
  .ZN(_1204_)
);

INV_X1 _5305_ (
  .A(\d_pipe[6][23] ),
  .ZN(_1205_)
);

NAND3_X1 _5306_ (
  .A1(_1202_),
  .A2(_1205_),
  .A3(_1154_),
  .ZN(_1206_)
);

NAND3_X1 _5307_ (
  .A1(_1204_),
  .A2(_1149_),
  .A3(_1206_),
  .ZN(_1207_)
);

OAI21_X1 _5308_ (
  .A(_1207_),
  .B1(_1149_),
  .B2(_0070_),
  .ZN(_4498_)
);

XNOR2_X1 _5309_ (
  .A(_4503_),
  .B(\d_pipe[5][14] ),
  .ZN(_1208_)
);

BUF_X1 _5310_ (
  .A(_0654_),
  .Z(_1209_)
);

NAND2_X1 _5311_ (
  .A1(_1208_),
  .A2(_1209_),
  .ZN(_1210_)
);

OAI21_X1 _5312_ (
  .A(_1210_),
  .B1(_1209_),
  .B2(_0071_),
  .ZN(_4507_)
);

INV_X2 _5313_ (
  .A(\d_pipe[5][14] ),
  .ZN(_1211_)
);

INV_X1 _5314_ (
  .A(\d_pipe[5][13] ),
  .ZN(_1212_)
);

NAND3_X2 _5315_ (
  .A1(_1211_),
  .A2(_1212_),
  .A3(_4501_),
  .ZN(_1213_)
);

INV_X1 _5316_ (
  .A(_1213_),
  .ZN(_1214_)
);

INV_X4 _5317_ (
  .A(\d_pipe[5][15] ),
  .ZN(_1215_)
);

OAI21_X1 _5318_ (
  .A(_0655_),
  .B1(_1214_),
  .B2(_1215_),
  .ZN(_1216_)
);

NAND2_X1 _5319_ (
  .A1(_1214_),
  .A2(_1215_),
  .ZN(_1217_)
);

INV_X1 _5320_ (
  .A(_1217_),
  .ZN(_1218_)
);

OAI22_X1 _5321_ (
  .A1(_1216_),
  .A2(_1218_),
  .B1(_0072_),
  .B2(_1209_),
  .ZN(_4510_)
);

NAND3_X2 _5322_ (
  .A1(_1211_),
  .A2(_1215_),
  .A3(_4503_),
  .ZN(_1219_)
);

BUF_X4 _5323_ (
  .A(\d_pipe[5][16] ),
  .Z(_1220_)
);

OR2_X1 _5324_ (
  .A1(_1219_),
  .A2(_1220_),
  .ZN(_1221_)
);

NAND2_X1 _5325_ (
  .A1(_1219_),
  .A2(_1220_),
  .ZN(_1222_)
);

NAND3_X1 _5326_ (
  .A1(_1221_),
  .A2(_0655_),
  .A3(_1222_),
  .ZN(_1223_)
);

OAI21_X1 _5327_ (
  .A(_1223_),
  .B1(_1209_),
  .B2(_0073_),
  .ZN(_4513_)
);

BUF_X4 _5328_ (
  .A(\d_pipe[5][17] ),
  .Z(_1224_)
);

INV_X2 _5329_ (
  .A(_1224_),
  .ZN(_1225_)
);

OAI21_X1 _5330_ (
  .A(_1225_),
  .B1(_1217_),
  .B2(_1220_),
  .ZN(_1226_)
);

INV_X1 _5331_ (
  .A(_1226_),
  .ZN(_1227_)
);

NOR3_X1 _5332_ (
  .A1(_1217_),
  .A2(_1220_),
  .A3(_1225_),
  .ZN(_1228_)
);

OAI21_X1 _5333_ (
  .A(_1209_),
  .B1(_1227_),
  .B2(_1228_),
  .ZN(_1229_)
);

OAI21_X1 _5334_ (
  .A(_1229_),
  .B1(_1209_),
  .B2(_0074_),
  .ZN(_4516_)
);

NOR2_X1 _5335_ (
  .A1(_1221_),
  .A2(_1224_),
  .ZN(_1230_)
);

INV_X1 _5336_ (
  .A(\d_pipe[5][18] ),
  .ZN(_1231_)
);

OAI21_X1 _5337_ (
  .A(_0655_),
  .B1(_1230_),
  .B2(_1231_),
  .ZN(_1232_)
);

NOR3_X1 _5338_ (
  .A1(_1221_),
  .A2(_1224_),
  .A3(\d_pipe[5][18] ),
  .ZN(_1233_)
);

OAI22_X1 _5339_ (
  .A1(_1232_),
  .A2(_1233_),
  .B1(_0075_),
  .B2(_1209_),
  .ZN(_4519_)
);

OR2_X1 _5340_ (
  .A1(_0655_),
  .A2(_0076_),
  .ZN(_1234_)
);

INV_X2 _5341_ (
  .A(_1220_),
  .ZN(_1235_)
);

NAND4_X1 _5342_ (
  .A1(_1225_),
  .A2(_1231_),
  .A3(_1215_),
  .A4(_1235_),
  .ZN(_1236_)
);

NOR2_X1 _5343_ (
  .A1(_1236_),
  .A2(_1213_),
  .ZN(_1237_)
);

INV_X1 _5344_ (
  .A(\d_pipe[5][19] ),
  .ZN(_1238_)
);

XNOR2_X1 _5345_ (
  .A(_1237_),
  .B(_1238_),
  .ZN(_1239_)
);

OAI21_X2 _5346_ (
  .A(_1234_),
  .B1(_1239_),
  .B2(\s_pipe[5][24] ),
  .ZN(_4522_)
);

OR2_X1 _5347_ (
  .A1(_0655_),
  .A2(_0077_),
  .ZN(_1240_)
);

NOR2_X4 _5348_ (
  .A1(_1220_),
  .A2(_1224_),
  .ZN(_1241_)
);

NOR2_X1 _5349_ (
  .A1(\d_pipe[5][18] ),
  .A2(\d_pipe[5][19] ),
  .ZN(_1242_)
);

NAND2_X2 _5350_ (
  .A1(_1241_),
  .A2(_1242_),
  .ZN(_1243_)
);

NOR2_X4 _5351_ (
  .A1(_1243_),
  .A2(_1219_),
  .ZN(_1244_)
);

INV_X1 _5352_ (
  .A(\d_pipe[5][20] ),
  .ZN(_1245_)
);

XNOR2_X1 _5353_ (
  .A(_1244_),
  .B(_1245_),
  .ZN(_1246_)
);

OAI21_X1 _5354_ (
  .A(_1240_),
  .B1(_1246_),
  .B2(\s_pipe[5][24] ),
  .ZN(_4525_)
);

NAND4_X1 _5355_ (
  .A1(_1215_),
  .A2(_1235_),
  .A3(_1211_),
  .A4(_1212_),
  .ZN(_1247_)
);

NAND2_X1 _5356_ (
  .A1(_1225_),
  .A2(_1231_),
  .ZN(_1248_)
);

NAND2_X1 _5357_ (
  .A1(_1238_),
  .A2(_1245_),
  .ZN(_1249_)
);

NOR3_X2 _5358_ (
  .A1(_1247_),
  .A2(_1248_),
  .A3(_1249_),
  .ZN(_1250_)
);

BUF_X4 _5359_ (
  .A(\d_pipe[5][21] ),
  .Z(_1251_)
);

NAND3_X1 _5360_ (
  .A1(_1250_),
  .A2(_4501_),
  .A3(_1251_),
  .ZN(_1252_)
);

INV_X1 _5361_ (
  .A(_1252_),
  .ZN(_1253_)
);

AOI21_X1 _5362_ (
  .A(_1251_),
  .B1(_1250_),
  .B2(_4501_),
  .ZN(_1254_)
);

OAI21_X1 _5363_ (
  .A(_1209_),
  .B1(_1253_),
  .B2(_1254_),
  .ZN(_1255_)
);

OR2_X1 _5364_ (
  .A1(_0655_),
  .A2(_0078_),
  .ZN(_1256_)
);

NAND2_X1 _5365_ (
  .A1(_1255_),
  .A2(_1256_),
  .ZN(_4528_)
);

INV_X1 _5366_ (
  .A(_1244_),
  .ZN(_1257_)
);

NOR2_X4 _5367_ (
  .A1(\d_pipe[5][20] ),
  .A2(_1251_),
  .ZN(_1258_)
);

INV_X1 _5368_ (
  .A(\d_pipe[5][22] ),
  .ZN(_1259_)
);

NAND2_X2 _5369_ (
  .A1(_1258_),
  .A2(_1259_),
  .ZN(_1260_)
);

OAI21_X1 _5370_ (
  .A(_0655_),
  .B1(_1257_),
  .B2(_1260_),
  .ZN(_1261_)
);

AOI21_X1 _5371_ (
  .A(_1259_),
  .B1(_1244_),
  .B2(_1258_),
  .ZN(_1262_)
);

OAI22_X1 _5372_ (
  .A1(_1261_),
  .A2(_1262_),
  .B1(_0079_),
  .B2(_1209_),
  .ZN(_4531_)
);

INV_X1 _5373_ (
  .A(_1251_),
  .ZN(_1263_)
);

NAND4_X1 _5374_ (
  .A1(_1263_),
  .A2(_1259_),
  .A3(_1238_),
  .A4(_1245_),
  .ZN(_1264_)
);

NOR2_X2 _5375_ (
  .A1(_1236_),
  .A2(_1264_),
  .ZN(_1265_)
);

INV_X1 _5376_ (
  .A(_1265_),
  .ZN(_1266_)
);

OAI21_X1 _5377_ (
  .A(\d_pipe[5][23] ),
  .B1(_1266_),
  .B2(_1213_),
  .ZN(_1267_)
);

INV_X1 _5378_ (
  .A(\d_pipe[5][23] ),
  .ZN(_1268_)
);

NAND3_X1 _5379_ (
  .A1(_1265_),
  .A2(_1268_),
  .A3(_1214_),
  .ZN(_1269_)
);

NAND3_X1 _5380_ (
  .A1(_1267_),
  .A2(_0655_),
  .A3(_1269_),
  .ZN(_1270_)
);

OAI21_X1 _5381_ (
  .A(_1270_),
  .B1(_1209_),
  .B2(_0080_),
  .ZN(_4534_)
);

XNOR2_X1 _5382_ (
  .A(_4539_),
  .B(\d_pipe[4][14] ),
  .ZN(_1271_)
);

BUF_X1 _5383_ (
  .A(_0657_),
  .Z(_1272_)
);

NAND2_X1 _5384_ (
  .A1(_1271_),
  .A2(_1272_),
  .ZN(_1273_)
);

OAI21_X1 _5385_ (
  .A(_1273_),
  .B1(_1272_),
  .B2(_0081_),
  .ZN(_4543_)
);

INV_X2 _5386_ (
  .A(\d_pipe[4][14] ),
  .ZN(_1274_)
);

INV_X1 _5387_ (
  .A(\d_pipe[4][13] ),
  .ZN(_1275_)
);

NAND3_X2 _5388_ (
  .A1(_1274_),
  .A2(_1275_),
  .A3(_4537_),
  .ZN(_1276_)
);

INV_X1 _5389_ (
  .A(_1276_),
  .ZN(_1277_)
);

INV_X4 _5390_ (
  .A(\d_pipe[4][15] ),
  .ZN(_1278_)
);

OAI21_X1 _5391_ (
  .A(_0658_),
  .B1(_1277_),
  .B2(_1278_),
  .ZN(_1279_)
);

NAND2_X1 _5392_ (
  .A1(_1277_),
  .A2(_1278_),
  .ZN(_1280_)
);

INV_X1 _5393_ (
  .A(_1280_),
  .ZN(_1281_)
);

OAI22_X1 _5394_ (
  .A1(_1279_),
  .A2(_1281_),
  .B1(_0082_),
  .B2(_1272_),
  .ZN(_4546_)
);

NAND3_X2 _5395_ (
  .A1(_1274_),
  .A2(_1278_),
  .A3(_4539_),
  .ZN(_1282_)
);

BUF_X4 _5396_ (
  .A(\d_pipe[4][16] ),
  .Z(_1283_)
);

OR2_X1 _5397_ (
  .A1(_1282_),
  .A2(_1283_),
  .ZN(_1284_)
);

NAND2_X1 _5398_ (
  .A1(_1282_),
  .A2(_1283_),
  .ZN(_1285_)
);

NAND3_X1 _5399_ (
  .A1(_1284_),
  .A2(_0658_),
  .A3(_1285_),
  .ZN(_1286_)
);

OAI21_X1 _5400_ (
  .A(_1286_),
  .B1(_1272_),
  .B2(_0083_),
  .ZN(_4549_)
);

BUF_X4 _5401_ (
  .A(\d_pipe[4][17] ),
  .Z(_1287_)
);

INV_X2 _5402_ (
  .A(_1287_),
  .ZN(_1288_)
);

OAI21_X1 _5403_ (
  .A(_1288_),
  .B1(_1280_),
  .B2(_1283_),
  .ZN(_1289_)
);

INV_X1 _5404_ (
  .A(_1289_),
  .ZN(_1290_)
);

NOR3_X1 _5405_ (
  .A1(_1280_),
  .A2(_1283_),
  .A3(_1288_),
  .ZN(_1291_)
);

OAI21_X1 _5406_ (
  .A(_1272_),
  .B1(_1290_),
  .B2(_1291_),
  .ZN(_1292_)
);

OAI21_X1 _5407_ (
  .A(_1292_),
  .B1(_1272_),
  .B2(_0084_),
  .ZN(_4552_)
);

NOR2_X1 _5408_ (
  .A1(_1284_),
  .A2(_1287_),
  .ZN(_1293_)
);

INV_X1 _5409_ (
  .A(\d_pipe[4][18] ),
  .ZN(_1294_)
);

OAI21_X1 _5410_ (
  .A(_0658_),
  .B1(_1293_),
  .B2(_1294_),
  .ZN(_1295_)
);

NOR3_X1 _5411_ (
  .A1(_1284_),
  .A2(_1287_),
  .A3(\d_pipe[4][18] ),
  .ZN(_1296_)
);

OAI22_X1 _5412_ (
  .A1(_1295_),
  .A2(_1296_),
  .B1(_0085_),
  .B2(_1272_),
  .ZN(_4555_)
);

OR2_X1 _5413_ (
  .A1(_0658_),
  .A2(_0086_),
  .ZN(_1297_)
);

INV_X2 _5414_ (
  .A(_1283_),
  .ZN(_1298_)
);

NAND4_X1 _5415_ (
  .A1(_1288_),
  .A2(_1294_),
  .A3(_1278_),
  .A4(_1298_),
  .ZN(_1299_)
);

NOR2_X1 _5416_ (
  .A1(_1299_),
  .A2(_1276_),
  .ZN(_1300_)
);

INV_X1 _5417_ (
  .A(\d_pipe[4][19] ),
  .ZN(_1301_)
);

XNOR2_X1 _5418_ (
  .A(_1300_),
  .B(_1301_),
  .ZN(_1302_)
);

OAI21_X1 _5419_ (
  .A(_1297_),
  .B1(_1302_),
  .B2(\s_pipe[4][24] ),
  .ZN(_4558_)
);

OR2_X1 _5420_ (
  .A1(_0658_),
  .A2(_0087_),
  .ZN(_1303_)
);

NOR2_X4 _5421_ (
  .A1(_1283_),
  .A2(_1287_),
  .ZN(_1304_)
);

NOR2_X1 _5422_ (
  .A1(\d_pipe[4][18] ),
  .A2(\d_pipe[4][19] ),
  .ZN(_1305_)
);

NAND2_X2 _5423_ (
  .A1(_1304_),
  .A2(_1305_),
  .ZN(_1306_)
);

NOR2_X4 _5424_ (
  .A1(_1306_),
  .A2(_1282_),
  .ZN(_1307_)
);

INV_X1 _5425_ (
  .A(\d_pipe[4][20] ),
  .ZN(_1308_)
);

XNOR2_X1 _5426_ (
  .A(_1307_),
  .B(_1308_),
  .ZN(_1309_)
);

OAI21_X1 _5427_ (
  .A(_1303_),
  .B1(_1309_),
  .B2(\s_pipe[4][24] ),
  .ZN(_4561_)
);

NAND4_X1 _5428_ (
  .A1(_1278_),
  .A2(_1298_),
  .A3(_1274_),
  .A4(_1275_),
  .ZN(_1310_)
);

NAND2_X1 _5429_ (
  .A1(_1288_),
  .A2(_1294_),
  .ZN(_1311_)
);

NAND2_X1 _5430_ (
  .A1(_1301_),
  .A2(_1308_),
  .ZN(_1312_)
);

NOR3_X2 _5431_ (
  .A1(_1310_),
  .A2(_1311_),
  .A3(_1312_),
  .ZN(_1313_)
);

BUF_X4 _5432_ (
  .A(\d_pipe[4][21] ),
  .Z(_1314_)
);

NAND3_X1 _5433_ (
  .A1(_1313_),
  .A2(_4537_),
  .A3(_1314_),
  .ZN(_1315_)
);

INV_X1 _5434_ (
  .A(_1315_),
  .ZN(_1316_)
);

AOI21_X1 _5435_ (
  .A(_1314_),
  .B1(_1313_),
  .B2(_4537_),
  .ZN(_1317_)
);

OAI21_X1 _5436_ (
  .A(_1272_),
  .B1(_1316_),
  .B2(_1317_),
  .ZN(_1318_)
);

OR2_X1 _5437_ (
  .A1(_0658_),
  .A2(_0088_),
  .ZN(_1319_)
);

NAND2_X1 _5438_ (
  .A1(_1318_),
  .A2(_1319_),
  .ZN(_4564_)
);

INV_X1 _5439_ (
  .A(_1307_),
  .ZN(_1320_)
);

NOR2_X4 _5440_ (
  .A1(\d_pipe[4][20] ),
  .A2(_1314_),
  .ZN(_1321_)
);

INV_X1 _5441_ (
  .A(\d_pipe[4][22] ),
  .ZN(_1322_)
);

NAND2_X2 _5442_ (
  .A1(_1321_),
  .A2(_1322_),
  .ZN(_1323_)
);

OAI21_X1 _5443_ (
  .A(_0658_),
  .B1(_1320_),
  .B2(_1323_),
  .ZN(_1324_)
);

AOI21_X1 _5444_ (
  .A(_1322_),
  .B1(_1307_),
  .B2(_1321_),
  .ZN(_1325_)
);

OAI22_X1 _5445_ (
  .A1(_1324_),
  .A2(_1325_),
  .B1(_0089_),
  .B2(_1272_),
  .ZN(_4567_)
);

INV_X1 _5446_ (
  .A(_1314_),
  .ZN(_1326_)
);

NAND4_X1 _5447_ (
  .A1(_1326_),
  .A2(_1322_),
  .A3(_1301_),
  .A4(_1308_),
  .ZN(_1327_)
);

NOR2_X1 _5448_ (
  .A1(_1299_),
  .A2(_1327_),
  .ZN(_1328_)
);

INV_X1 _5449_ (
  .A(_1328_),
  .ZN(_1329_)
);

OAI21_X1 _5450_ (
  .A(\d_pipe[4][23] ),
  .B1(_1329_),
  .B2(_1276_),
  .ZN(_1330_)
);

INV_X1 _5451_ (
  .A(\d_pipe[4][23] ),
  .ZN(_1331_)
);

NAND3_X1 _5452_ (
  .A1(_1328_),
  .A2(_1331_),
  .A3(_1277_),
  .ZN(_1332_)
);

NAND3_X1 _5453_ (
  .A1(_1330_),
  .A2(_0658_),
  .A3(_1332_),
  .ZN(_1333_)
);

OAI21_X1 _5454_ (
  .A(_1333_),
  .B1(_1272_),
  .B2(_0090_),
  .ZN(_4570_)
);

INV_X1 _5455_ (
  .A(d[11]),
  .ZN(_4282_)
);

INV_X1 _5456_ (
  .A(d[10]),
  .ZN(_4279_)
);

INV_X1 _5457_ (
  .A(d[4]),
  .ZN(_4261_)
);

INV_X1 _5458_ (
  .A(d[3]),
  .ZN(_4258_)
);

INV_X1 _5459_ (
  .A(d[1]),
  .ZN(_4252_)
);

BUF_X2 _5460_ (
  .A(ena),
  .Z(_1334_)
);

BUF_X2 _5461_ (
  .A(_1334_),
  .Z(_1335_)
);

BUF_X2 _5462_ (
  .A(_1335_),
  .Z(_1336_)
);

INV_X2 _5464_ (
  .A(_1334_),
  .ZN(_1337_)
);

BUF_X1 _5465_ (
  .A(_1337_),
  .Z(_1338_)
);

BUF_X4 _5467_ (
  .A(_1337_),
  .Z(_1340_)
);

BUF_X2 _5468_ (
  .A(_1340_),
  .Z(_1341_)
);

INV_X1 _5470_ (
  .A(_4069_),
  .ZN(_1342_)
);

NAND2_X1 _5471_ (
  .A1(_1342_),
  .A2(_4293_),
  .ZN(_1343_)
);

BUF_X4 _5474_ (
  .A(_1334_),
  .Z(_1346_)
);

BUF_X8 _5475_ (
  .A(_1346_),
  .Z(_1347_)
);

BUF_X2 _5476_ (
  .A(_1347_),
  .Z(_1348_)
);

BUF_X2 _5478_ (
  .A(_1346_),
  .Z(_1350_)
);

BUF_X2 _5479_ (
  .A(_1350_),
  .Z(_1351_)
);

BUF_X4 _5482_ (
  .A(_1347_),
  .Z(_1353_)
);

INV_X1 _5490_ (
  .A(_4296_),
  .ZN(_1361_)
);

BUF_X2 _5492_ (
  .A(_1350_),
  .Z(_1363_)
);

BUF_X4 _5494_ (
  .A(_1347_),
  .Z(_1364_)
);

NOR2_X1 _5496_ (
  .A1(_4292_),
  .A2(_4295_),
  .ZN(_1366_)
);

INV_X1 _5497_ (
  .A(_4295_),
  .ZN(_1367_)
);

AOI22_X2 _5498_ (
  .A1(_1366_),
  .A2(_1343_),
  .B1(_1367_),
  .B2(_1361_),
  .ZN(_1368_)
);

BUF_X4 _5499_ (
  .A(_4299_),
  .Z(_1369_)
);

BUF_X4 _5502_ (
  .A(_1347_),
  .Z(_1371_)
);

INV_X1 _5504_ (
  .A(_4298_),
  .ZN(_1373_)
);

BUF_X4 _5510_ (
  .A(_4302_),
  .Z(_1379_)
);

BUF_X2 _5512_ (
  .A(_1350_),
  .Z(_1381_)
);

INV_X1 _5515_ (
  .A(_4301_),
  .ZN(_1383_)
);

INV_X1 _5516_ (
  .A(_1379_),
  .ZN(_1384_)
);

OAI21_X2 _5517_ (
  .A(_1383_),
  .B1(_1384_),
  .B2(_1373_),
  .ZN(_1385_)
);

NAND2_X1 _5518_ (
  .A1(_1369_),
  .A2(_1379_),
  .ZN(_1386_)
);

INV_X1 _5530_ (
  .A(_4304_),
  .ZN(_1397_)
);

INV_X1 _5537_ (
  .A(_4308_),
  .ZN(_1404_)
);

BUF_X4 _5539_ (
  .A(_1347_),
  .Z(_1406_)
);

BUF_X2 _5541_ (
  .A(_1350_),
  .Z(_1408_)
);

NAND2_X1 _5544_ (
  .A1(_4305_),
  .A2(_4308_),
  .ZN(_1410_)
);

NOR2_X2 _5545_ (
  .A1(_1386_),
  .A2(_1410_),
  .ZN(_1411_)
);

INV_X1 _5547_ (
  .A(_1410_),
  .ZN(_1413_)
);

NAND2_X1 _5548_ (
  .A1(_1385_),
  .A2(_1413_),
  .ZN(_1414_)
);

INV_X1 _5549_ (
  .A(_4307_),
  .ZN(_1415_)
);

OAI21_X1 _5550_ (
  .A(_1415_),
  .B1(_1404_),
  .B2(_1397_),
  .ZN(_1416_)
);

INV_X1 _5551_ (
  .A(_1416_),
  .ZN(_1417_)
);

NAND2_X1 _5552_ (
  .A1(_1414_),
  .A2(_1417_),
  .ZN(_1418_)
);

BUF_X2 _5560_ (
  .A(_1346_),
  .Z(_1426_)
);

BUF_X2 _5561_ (
  .A(_1426_),
  .Z(_1427_)
);

INV_X1 _5570_ (
  .A(_4310_),
  .ZN(_1435_)
);

INV_X1 _5579_ (
  .A(_4314_),
  .ZN(_1444_)
);

BUF_X4 _5581_ (
  .A(_1346_),
  .Z(_1446_)
);

BUF_X2 _5582_ (
  .A(_1446_),
  .Z(_1447_)
);

CLKBUF_X2 _5584_ (
  .A(_1340_),
  .Z(_1449_)
);

NAND2_X2 _5591_ (
  .A1(_4311_),
  .A2(_4314_),
  .ZN(_1455_)
);

INV_X2 _5594_ (
  .A(_1455_),
  .ZN(_1458_)
);

INV_X1 _5596_ (
  .A(_4313_),
  .ZN(_1460_)
);

OAI21_X1 _5597_ (
  .A(_1460_),
  .B1(_1444_),
  .B2(_1435_),
  .ZN(_1461_)
);

INV_X1 _5614_ (
  .A(_4316_),
  .ZN(_1477_)
);

INV_X1 _5622_ (
  .A(_4320_),
  .ZN(_1485_)
);

CLKBUF_X2 _5627_ (
  .A(_1340_),
  .Z(_1490_)
);

NAND2_X1 _5630_ (
  .A1(_4317_),
  .A2(_4320_),
  .ZN(_1492_)
);

INV_X1 _5631_ (
  .A(_1492_),
  .ZN(_1493_)
);

NAND2_X1 _5632_ (
  .A1(_1458_),
  .A2(_1493_),
  .ZN(_1494_)
);

INV_X2 _5633_ (
  .A(_1494_),
  .ZN(_1495_)
);

NAND2_X1 _5634_ (
  .A1(_1418_),
  .A2(_1495_),
  .ZN(_1496_)
);

AND2_X2 _5635_ (
  .A1(_1495_),
  .A2(_1411_),
  .ZN(_1497_)
);

NAND2_X1 _5636_ (
  .A1(_1368_),
  .A2(_1497_),
  .ZN(_1498_)
);

NAND2_X1 _5637_ (
  .A1(_1461_),
  .A2(_1493_),
  .ZN(_1499_)
);

INV_X1 _5638_ (
  .A(_4319_),
  .ZN(_1500_)
);

OAI21_X1 _5639_ (
  .A(_1500_),
  .B1(_1485_),
  .B2(_1477_),
  .ZN(_1501_)
);

INV_X1 _5640_ (
  .A(_1501_),
  .ZN(_1502_)
);

NAND2_X1 _5641_ (
  .A1(_1499_),
  .A2(_1502_),
  .ZN(_1503_)
);

INV_X1 _5642_ (
  .A(_1503_),
  .ZN(_1504_)
);

NAND3_X2 _5643_ (
  .A1(_1496_),
  .A2(_1498_),
  .A3(_1504_),
  .ZN(_1505_)
);

INV_X1 _5644_ (
  .A(_1505_),
  .ZN(_1506_)
);

NOR2_X2 _5645_ (
  .A1(_0904_),
  .A2(\d_pipe[11][23] ),
  .ZN(_1507_)
);

NAND2_X4 _5646_ (
  .A1(_0888_),
  .A2(_1507_),
  .ZN(_1508_)
);

NAND2_X2 _5647_ (
  .A1(_1508_),
  .A2(_0635_),
  .ZN(_1509_)
);

INV_X1 _5648_ (
  .A(\s_pipe[11][23] ),
  .ZN(_1510_)
);

NAND2_X1 _5649_ (
  .A1(_1509_),
  .A2(_1510_),
  .ZN(_1511_)
);

NAND3_X1 _5650_ (
  .A1(_1508_),
  .A2(_0635_),
  .A3(\s_pipe[11][23] ),
  .ZN(_1512_)
);

NAND2_X1 _5651_ (
  .A1(_1511_),
  .A2(_1512_),
  .ZN(_1513_)
);

NAND2_X1 _5652_ (
  .A1(_1506_),
  .A2(_1513_),
  .ZN(_1514_)
);

NAND2_X1 _5653_ (
  .A1(_1509_),
  .A2(\s_pipe[11][23] ),
  .ZN(_1515_)
);

NAND3_X1 _5654_ (
  .A1(_1508_),
  .A2(_0635_),
  .A3(_1510_),
  .ZN(_1516_)
);

NAND2_X1 _5655_ (
  .A1(_1515_),
  .A2(_1516_),
  .ZN(_1517_)
);

NAND2_X1 _5656_ (
  .A1(_1517_),
  .A2(_1505_),
  .ZN(_1518_)
);

NAND3_X1 _5657_ (
  .A1(_1514_),
  .A2(_1518_),
  .A3(_1447_),
  .ZN(_1519_)
);

BUF_X1 _5658_ (
  .A(\s_pipe[12][24] ),
  .Z(_1520_)
);

NAND2_X1 _5659_ (
  .A1(_1490_),
  .A2(_1520_),
  .ZN(_1521_)
);

NAND2_X1 _5660_ (
  .A1(_1519_),
  .A2(_1521_),
  .ZN(_0156_)
);

BUF_X2 _5661_ (
  .A(_1337_),
  .Z(_1522_)
);

NAND2_X1 _5662_ (
  .A1(_1522_),
  .A2(\d_pipe[3][12] ),
  .ZN(_1523_)
);

BUF_X2 _5663_ (
  .A(_1522_),
  .Z(_1524_)
);

INV_X1 _5664_ (
  .A(\d_pipe[2][12] ),
  .ZN(_1525_)
);

OAI21_X1 _5665_ (
  .A(_1523_),
  .B1(_1524_),
  .B2(_1525_),
  .ZN(_0157_)
);

BUF_X4 _5666_ (
  .A(_1346_),
  .Z(_1526_)
);

BUF_X2 _5667_ (
  .A(_1526_),
  .Z(_1527_)
);

NAND2_X1 _5668_ (
  .A1(\d_pipe[2][13] ),
  .A2(_1527_),
  .ZN(_1528_)
);

BUF_X2 _5669_ (
  .A(_1426_),
  .Z(_1529_)
);

OAI21_X1 _5670_ (
  .A(_1528_),
  .B1(_0748_),
  .B2(_1529_),
  .ZN(_0158_)
);

NAND2_X1 _5671_ (
  .A1(\d_pipe[2][14] ),
  .A2(_1527_),
  .ZN(_1530_)
);

BUF_X2 _5672_ (
  .A(_1426_),
  .Z(_1531_)
);

OAI21_X1 _5673_ (
  .A(_1530_),
  .B1(_0747_),
  .B2(_1531_),
  .ZN(_0159_)
);

NAND2_X1 _5674_ (
  .A1(\d_pipe[2][15] ),
  .A2(_1527_),
  .ZN(_1532_)
);

BUF_X2 _5675_ (
  .A(_1426_),
  .Z(_1533_)
);

OAI21_X1 _5676_ (
  .A(_1532_),
  .B1(_0751_),
  .B2(_1533_),
  .ZN(_0160_)
);

NAND2_X1 _5677_ (
  .A1(_0690_),
  .A2(_1527_),
  .ZN(_1534_)
);

BUF_X2 _5678_ (
  .A(_1426_),
  .Z(_1535_)
);

OAI21_X1 _5679_ (
  .A(_1534_),
  .B1(_0760_),
  .B2(_1535_),
  .ZN(_0161_)
);

NAND2_X1 _5680_ (
  .A1(_0695_),
  .A2(_1527_),
  .ZN(_1536_)
);

OAI21_X1 _5681_ (
  .A(_1536_),
  .B1(_0764_),
  .B2(_1535_),
  .ZN(_0162_)
);

BUF_X2 _5682_ (
  .A(_1526_),
  .Z(_1537_)
);

NAND2_X1 _5683_ (
  .A1(_0701_),
  .A2(_1537_),
  .ZN(_1538_)
);

BUF_X2 _5684_ (
  .A(_1426_),
  .Z(_1539_)
);

OAI21_X1 _5685_ (
  .A(_1538_),
  .B1(_0768_),
  .B2(_1539_),
  .ZN(_0163_)
);

NAND2_X1 _5686_ (
  .A1(\d_pipe[2][19] ),
  .A2(_1537_),
  .ZN(_1540_)
);

OAI21_X1 _5687_ (
  .A(_1540_),
  .B1(_0784_),
  .B2(_1539_),
  .ZN(_0164_)
);

NAND2_X1 _5688_ (
  .A1(\d_pipe[2][20] ),
  .A2(_1537_),
  .ZN(_1541_)
);

OAI21_X1 _5689_ (
  .A(_1541_),
  .B1(_0780_),
  .B2(_1539_),
  .ZN(_0165_)
);

NAND2_X1 _5690_ (
  .A1(_0722_),
  .A2(_1537_),
  .ZN(_1542_)
);

OAI21_X1 _5691_ (
  .A(_1542_),
  .B1(_0789_),
  .B2(_1539_),
  .ZN(_0166_)
);

NAND2_X1 _5692_ (
  .A1(\d_pipe[2][22] ),
  .A2(_1537_),
  .ZN(_1543_)
);

OAI21_X1 _5693_ (
  .A(_1543_),
  .B1(_0794_),
  .B2(_1539_),
  .ZN(_0167_)
);

BUF_X2 _5694_ (
  .A(_1526_),
  .Z(_1544_)
);

NAND2_X1 _5695_ (
  .A1(_0738_),
  .A2(_1544_),
  .ZN(_1545_)
);

OAI21_X1 _5696_ (
  .A(_1545_),
  .B1(_0802_),
  .B2(_1539_),
  .ZN(_0168_)
);

BUF_X2 _5697_ (
  .A(_1446_),
  .Z(_1546_)
);

NAND2_X1 _5698_ (
  .A1(_1546_),
  .A2(\d_pipe[1][12] ),
  .ZN(_1547_)
);

BUF_X2 _5699_ (
  .A(_1350_),
  .Z(_1548_)
);

OAI21_X1 _5700_ (
  .A(_1547_),
  .B1(_1548_),
  .B2(_1525_),
  .ZN(_0169_)
);

NAND2_X1 _5701_ (
  .A1(\d_pipe[1][13] ),
  .A2(_1544_),
  .ZN(_1549_)
);

OAI21_X1 _5702_ (
  .A(_1549_),
  .B1(_0660_),
  .B2(_1539_),
  .ZN(_0170_)
);

NAND2_X1 _5703_ (
  .A1(\d_pipe[1][14] ),
  .A2(_1544_),
  .ZN(_1550_)
);

OAI21_X1 _5704_ (
  .A(_1550_),
  .B1(_0661_),
  .B2(_1539_),
  .ZN(_0171_)
);

NAND2_X1 _5705_ (
  .A1(\d_pipe[1][15] ),
  .A2(_1544_),
  .ZN(_1551_)
);

BUF_X2 _5706_ (
  .A(_1426_),
  .Z(_1552_)
);

OAI21_X1 _5707_ (
  .A(_1551_),
  .B1(_0663_),
  .B2(_1552_),
  .ZN(_0172_)
);

NAND2_X1 _5708_ (
  .A1(_0806_),
  .A2(_1544_),
  .ZN(_1553_)
);

OAI21_X1 _5709_ (
  .A(_1553_),
  .B1(_0717_),
  .B2(_1552_),
  .ZN(_0173_)
);

NAND2_X1 _5710_ (
  .A1(_0811_),
  .A2(_1544_),
  .ZN(_1554_)
);

OAI21_X1 _5711_ (
  .A(_1554_),
  .B1(_0696_),
  .B2(_1552_),
  .ZN(_0174_)
);

NAND2_X1 _5712_ (
  .A1(\d_pipe[1][18] ),
  .A2(_1544_),
  .ZN(_1555_)
);

OAI21_X1 _5713_ (
  .A(_1555_),
  .B1(_0702_),
  .B2(_1552_),
  .ZN(_0175_)
);

NAND2_X1 _5714_ (
  .A1(\d_pipe[1][19] ),
  .A2(_1544_),
  .ZN(_1556_)
);

OAI21_X1 _5715_ (
  .A(_1556_),
  .B1(_0706_),
  .B2(_1552_),
  .ZN(_0176_)
);

NAND2_X1 _5716_ (
  .A1(\d_pipe[1][20] ),
  .A2(_1544_),
  .ZN(_1557_)
);

OAI21_X1 _5717_ (
  .A(_1557_),
  .B1(_0715_),
  .B2(_1552_),
  .ZN(_0177_)
);

BUF_X2 _5718_ (
  .A(_1526_),
  .Z(_1558_)
);

NAND2_X1 _5719_ (
  .A1(\d_pipe[1][21] ),
  .A2(_1558_),
  .ZN(_1559_)
);

OAI21_X1 _5720_ (
  .A(_1559_),
  .B1(_0735_),
  .B2(_1552_),
  .ZN(_0178_)
);

NAND2_X1 _5721_ (
  .A1(\d_pipe[1][22] ),
  .A2(_1558_),
  .ZN(_1560_)
);

OAI21_X1 _5722_ (
  .A(_1560_),
  .B1(_0730_),
  .B2(_1531_),
  .ZN(_0179_)
);

NAND2_X1 _5723_ (
  .A1(_1522_),
  .A2(_0738_),
  .ZN(_1561_)
);

BUF_X2 _5724_ (
  .A(_1340_),
  .Z(_1562_)
);

OAI21_X1 _5725_ (
  .A(_1561_),
  .B1(_0851_),
  .B2(_1562_),
  .ZN(_0180_)
);

BUF_X2 _5726_ (
  .A(_1335_),
  .Z(_1563_)
);

MUX2_X1 _5727_ (
  .A(\s_pipe[1][1] ),
  .B(z[0]),
  .S(_1563_),
  .Z(_0181_)
);

MUX2_X1 _5728_ (
  .A(\s_pipe[1][2] ),
  .B(z[1]),
  .S(_1563_),
  .Z(_0182_)
);

BUF_X2 _5729_ (
  .A(_1346_),
  .Z(_1564_)
);

MUX2_X1 _5730_ (
  .A(\s_pipe[1][3] ),
  .B(z[2]),
  .S(_1564_),
  .Z(_0183_)
);

MUX2_X1 _5731_ (
  .A(\s_pipe[1][4] ),
  .B(z[3]),
  .S(_1564_),
  .Z(_0184_)
);

MUX2_X1 _5732_ (
  .A(\s_pipe[1][5] ),
  .B(z[4]),
  .S(_1564_),
  .Z(_0185_)
);

MUX2_X1 _5733_ (
  .A(\s_pipe[1][6] ),
  .B(z[5]),
  .S(_1564_),
  .Z(_0186_)
);

MUX2_X1 _5734_ (
  .A(\s_pipe[1][7] ),
  .B(z[6]),
  .S(_1564_),
  .Z(_0187_)
);

BUF_X2 _5735_ (
  .A(_1346_),
  .Z(_1565_)
);

MUX2_X1 _5736_ (
  .A(\s_pipe[1][8] ),
  .B(z[7]),
  .S(_1565_),
  .Z(_0188_)
);

BUF_X2 _5737_ (
  .A(_1335_),
  .Z(_1566_)
);

MUX2_X1 _5738_ (
  .A(\s_pipe[1][9] ),
  .B(z[8]),
  .S(_1566_),
  .Z(_0189_)
);

MUX2_X1 _5739_ (
  .A(\s_pipe[1][10] ),
  .B(z[9]),
  .S(_1565_),
  .Z(_0190_)
);

MUX2_X1 _5740_ (
  .A(\s_pipe[1][11] ),
  .B(z[10]),
  .S(_1565_),
  .Z(_0191_)
);

NAND2_X1 _5741_ (
  .A1(_1522_),
  .A2(\s_pipe[1][12] ),
  .ZN(_1567_)
);

OAI21_X1 _5742_ (
  .A(_1567_),
  .B1(_4123_),
  .B2(_1341_),
  .ZN(_0192_)
);

MUX2_X1 _5743_ (
  .A(\s_pipe[1][13] ),
  .B(_0143_),
  .S(_1565_),
  .Z(_0193_)
);

INV_X1 _5744_ (
  .A(_4257_),
  .ZN(_1568_)
);

NAND2_X1 _5745_ (
  .A1(_1568_),
  .A2(_4065_),
  .ZN(_1569_)
);

INV_X1 _5746_ (
  .A(_4065_),
  .ZN(_1570_)
);

NAND2_X1 _5747_ (
  .A1(_1570_),
  .A2(_4257_),
  .ZN(_1571_)
);

BUF_X2 _5748_ (
  .A(_1347_),
  .Z(_1572_)
);

NAND3_X1 _5749_ (
  .A1(_1569_),
  .A2(_1571_),
  .A3(_1572_),
  .ZN(_1573_)
);

INV_X1 _5750_ (
  .A(\s_pipe[1][14] ),
  .ZN(_1574_)
);

OAI21_X1 _5751_ (
  .A(_1573_),
  .B1(_1351_),
  .B2(_1574_),
  .ZN(_0194_)
);

NOR2_X1 _5752_ (
  .A1(_1371_),
  .A2(\s_pipe[1][15] ),
  .ZN(_1575_)
);

INV_X1 _5753_ (
  .A(_4256_),
  .ZN(_1576_)
);

INV_X1 _5754_ (
  .A(_4253_),
  .ZN(_1577_)
);

OAI21_X2 _5755_ (
  .A(_1576_),
  .B1(_1568_),
  .B2(_1577_),
  .ZN(_1578_)
);

INV_X1 _5756_ (
  .A(_1578_),
  .ZN(_1579_)
);

NAND2_X1 _5757_ (
  .A1(_4254_),
  .A2(_4257_),
  .ZN(_1580_)
);

INV_X1 _5758_ (
  .A(_1580_),
  .ZN(_1581_)
);

INV_X1 _5759_ (
  .A(_4064_),
  .ZN(_1582_)
);

NAND2_X1 _5760_ (
  .A1(_1581_),
  .A2(_1582_),
  .ZN(_1583_)
);

NAND2_X2 _5761_ (
  .A1(_1579_),
  .A2(_1583_),
  .ZN(_1584_)
);

BUF_X2 _5762_ (
  .A(_4260_),
  .Z(_1585_)
);

XNOR2_X1 _5763_ (
  .A(_1584_),
  .B(_1585_),
  .ZN(_1586_)
);

BUF_X2 _5764_ (
  .A(_1350_),
  .Z(_1587_)
);

AOI21_X1 _5765_ (
  .A(_1575_),
  .B1(_1586_),
  .B2(_1587_),
  .ZN(_0195_)
);

NOR2_X1 _5766_ (
  .A1(_1364_),
  .A2(\s_pipe[1][16] ),
  .ZN(_1588_)
);

INV_X1 _5767_ (
  .A(_4259_),
  .ZN(_1589_)
);

INV_X1 _5768_ (
  .A(_1585_),
  .ZN(_1590_)
);

OAI21_X2 _5769_ (
  .A(_1589_),
  .B1(_1590_),
  .B2(_1576_),
  .ZN(_1591_)
);

INV_X1 _5770_ (
  .A(_1591_),
  .ZN(_1592_)
);

NAND2_X1 _5771_ (
  .A1(_4257_),
  .A2(_1585_),
  .ZN(_1593_)
);

INV_X1 _5772_ (
  .A(_1593_),
  .ZN(_1594_)
);

NAND2_X1 _5773_ (
  .A1(_1594_),
  .A2(_1570_),
  .ZN(_1595_)
);

NAND2_X2 _5774_ (
  .A1(_1592_),
  .A2(_1595_),
  .ZN(_1596_)
);

BUF_X2 _5775_ (
  .A(_4263_),
  .Z(_1597_)
);

XNOR2_X1 _5776_ (
  .A(_1596_),
  .B(_1597_),
  .ZN(_1598_)
);

AOI21_X1 _5777_ (
  .A(_1588_),
  .B1(_1598_),
  .B2(_1381_),
  .ZN(_0196_)
);

INV_X1 _5778_ (
  .A(_4262_),
  .ZN(_1599_)
);

INV_X1 _5779_ (
  .A(_1597_),
  .ZN(_1600_)
);

OAI21_X2 _5780_ (
  .A(_1599_),
  .B1(_1600_),
  .B2(_1589_),
  .ZN(_1601_)
);

NAND2_X1 _5781_ (
  .A1(_1585_),
  .A2(_1597_),
  .ZN(_1602_)
);

INV_X2 _5782_ (
  .A(_1602_),
  .ZN(_1603_)
);

AOI21_X1 _5783_ (
  .A(_1601_),
  .B1(_1584_),
  .B2(_1603_),
  .ZN(_1604_)
);

INV_X1 _5784_ (
  .A(_4266_),
  .ZN(_1605_)
);

OR2_X1 _5785_ (
  .A1(_1604_),
  .A2(_1605_),
  .ZN(_1606_)
);

NAND2_X1 _5786_ (
  .A1(_1604_),
  .A2(_1605_),
  .ZN(_1607_)
);

NAND3_X1 _5787_ (
  .A1(_1606_),
  .A2(_1406_),
  .A3(_1607_),
  .ZN(_1608_)
);

INV_X1 _5788_ (
  .A(\s_pipe[1][17] ),
  .ZN(_1609_)
);

OAI21_X1 _5789_ (
  .A(_1608_),
  .B1(_1351_),
  .B2(_1609_),
  .ZN(_0197_)
);

INV_X1 _5790_ (
  .A(_4265_),
  .ZN(_1610_)
);

OAI21_X2 _5791_ (
  .A(_1610_),
  .B1(_1605_),
  .B2(_1599_),
  .ZN(_1611_)
);

NAND2_X1 _5792_ (
  .A1(_1597_),
  .A2(_4266_),
  .ZN(_1612_)
);

INV_X2 _5793_ (
  .A(_1612_),
  .ZN(_1613_)
);

AOI21_X2 _5794_ (
  .A(_1611_),
  .B1(_1596_),
  .B2(_1613_),
  .ZN(_1614_)
);

INV_X1 _5795_ (
  .A(_4269_),
  .ZN(_1615_)
);

OR2_X2 _5796_ (
  .A1(_1614_),
  .A2(_1615_),
  .ZN(_1616_)
);

NAND2_X1 _5797_ (
  .A1(_1614_),
  .A2(_1615_),
  .ZN(_1617_)
);

NAND3_X1 _5798_ (
  .A1(_1616_),
  .A2(_1406_),
  .A3(_1617_),
  .ZN(_1618_)
);

INV_X1 _5799_ (
  .A(\s_pipe[1][18] ),
  .ZN(_1619_)
);

OAI21_X1 _5800_ (
  .A(_1618_),
  .B1(_1351_),
  .B2(_1619_),
  .ZN(_0198_)
);

NAND2_X1 _5801_ (
  .A1(_4266_),
  .A2(_4269_),
  .ZN(_1620_)
);

INV_X1 _5802_ (
  .A(_1620_),
  .ZN(_1621_)
);

NAND3_X1 _5803_ (
  .A1(_1584_),
  .A2(_1603_),
  .A3(_1621_),
  .ZN(_1622_)
);

NAND2_X1 _5804_ (
  .A1(_1601_),
  .A2(_1621_),
  .ZN(_1623_)
);

INV_X1 _5805_ (
  .A(_4268_),
  .ZN(_1624_)
);

OAI21_X1 _5806_ (
  .A(_1624_),
  .B1(_1615_),
  .B2(_1610_),
  .ZN(_1625_)
);

INV_X1 _5807_ (
  .A(_1625_),
  .ZN(_1626_)
);

NAND2_X1 _5808_ (
  .A1(_1623_),
  .A2(_1626_),
  .ZN(_1627_)
);

INV_X1 _5809_ (
  .A(_1627_),
  .ZN(_1628_)
);

NAND2_X1 _5810_ (
  .A1(_1622_),
  .A2(_1628_),
  .ZN(_1629_)
);

NAND2_X1 _5811_ (
  .A1(_1629_),
  .A2(_4272_),
  .ZN(_1630_)
);

INV_X1 _5812_ (
  .A(_4272_),
  .ZN(_1631_)
);

NAND3_X1 _5813_ (
  .A1(_1622_),
  .A2(_1631_),
  .A3(_1628_),
  .ZN(_1632_)
);

NAND3_X1 _5814_ (
  .A1(_1630_),
  .A2(_1632_),
  .A3(_1348_),
  .ZN(_1633_)
);

BUF_X2 _5815_ (
  .A(_1350_),
  .Z(_1634_)
);

INV_X1 _5816_ (
  .A(\s_pipe[1][19] ),
  .ZN(_1635_)
);

OAI21_X1 _5817_ (
  .A(_1633_),
  .B1(_1634_),
  .B2(_1635_),
  .ZN(_0199_)
);

NAND2_X1 _5818_ (
  .A1(_4269_),
  .A2(_4272_),
  .ZN(_1636_)
);

INV_X1 _5819_ (
  .A(_1636_),
  .ZN(_1637_)
);

NAND3_X1 _5820_ (
  .A1(_1596_),
  .A2(_1613_),
  .A3(_1637_),
  .ZN(_1638_)
);

NAND2_X1 _5821_ (
  .A1(_1611_),
  .A2(_1637_),
  .ZN(_1639_)
);

INV_X1 _5822_ (
  .A(_4271_),
  .ZN(_1640_)
);

OAI21_X1 _5823_ (
  .A(_1640_),
  .B1(_1631_),
  .B2(_1624_),
  .ZN(_1641_)
);

INV_X1 _5824_ (
  .A(_1641_),
  .ZN(_1642_)
);

NAND2_X1 _5825_ (
  .A1(_1639_),
  .A2(_1642_),
  .ZN(_1643_)
);

INV_X1 _5826_ (
  .A(_1643_),
  .ZN(_1644_)
);

NAND2_X1 _5827_ (
  .A1(_1638_),
  .A2(_1644_),
  .ZN(_1645_)
);

NAND2_X1 _5828_ (
  .A1(_1645_),
  .A2(_4275_),
  .ZN(_1646_)
);

INV_X1 _5829_ (
  .A(_4275_),
  .ZN(_1647_)
);

NAND3_X1 _5830_ (
  .A1(_1638_),
  .A2(_1647_),
  .A3(_1644_),
  .ZN(_1648_)
);

NAND3_X1 _5831_ (
  .A1(_1646_),
  .A2(_1648_),
  .A3(_1348_),
  .ZN(_1649_)
);

INV_X1 _5832_ (
  .A(\s_pipe[1][20] ),
  .ZN(_1650_)
);

OAI21_X1 _5833_ (
  .A(_1649_),
  .B1(_1634_),
  .B2(_1650_),
  .ZN(_0200_)
);

NAND2_X1 _5834_ (
  .A1(_1578_),
  .A2(_1603_),
  .ZN(_1651_)
);

INV_X1 _5835_ (
  .A(_1601_),
  .ZN(_1652_)
);

NAND2_X1 _5836_ (
  .A1(_1651_),
  .A2(_1652_),
  .ZN(_1653_)
);

NAND2_X1 _5837_ (
  .A1(_4272_),
  .A2(_4275_),
  .ZN(_1654_)
);

NOR2_X1 _5838_ (
  .A1(_1620_),
  .A2(_1654_),
  .ZN(_1655_)
);

NAND2_X1 _5839_ (
  .A1(_1653_),
  .A2(_1655_),
  .ZN(_1656_)
);

INV_X1 _5840_ (
  .A(_1654_),
  .ZN(_1657_)
);

NAND2_X1 _5841_ (
  .A1(_1625_),
  .A2(_1657_),
  .ZN(_1658_)
);

INV_X1 _5842_ (
  .A(_4274_),
  .ZN(_1659_)
);

OAI21_X1 _5843_ (
  .A(_1659_),
  .B1(_1647_),
  .B2(_1640_),
  .ZN(_1660_)
);

INV_X1 _5844_ (
  .A(_1660_),
  .ZN(_1661_)
);

NAND2_X1 _5845_ (
  .A1(_1658_),
  .A2(_1661_),
  .ZN(_1662_)
);

INV_X1 _5846_ (
  .A(_1662_),
  .ZN(_1663_)
);

NAND4_X1 _5847_ (
  .A1(_1655_),
  .A2(_1603_),
  .A3(_1581_),
  .A4(_1582_),
  .ZN(_1664_)
);

NAND3_X1 _5848_ (
  .A1(_1656_),
  .A2(_1663_),
  .A3(_1664_),
  .ZN(_1665_)
);

NAND2_X1 _5849_ (
  .A1(_1665_),
  .A2(_4278_),
  .ZN(_1666_)
);

INV_X1 _5850_ (
  .A(_4278_),
  .ZN(_1667_)
);

NAND4_X1 _5851_ (
  .A1(_1656_),
  .A2(_1664_),
  .A3(_1663_),
  .A4(_1667_),
  .ZN(_1668_)
);

BUF_X2 _5852_ (
  .A(_1446_),
  .Z(_1669_)
);

NAND3_X1 _5853_ (
  .A1(_1666_),
  .A2(_1668_),
  .A3(_1669_),
  .ZN(_1670_)
);

NAND2_X1 _5854_ (
  .A1(_1490_),
  .A2(\s_pipe[1][21] ),
  .ZN(_1671_)
);

NAND2_X1 _5855_ (
  .A1(_1670_),
  .A2(_1671_),
  .ZN(_0201_)
);

NAND2_X1 _5856_ (
  .A1(_1591_),
  .A2(_1613_),
  .ZN(_1672_)
);

INV_X1 _5857_ (
  .A(_1611_),
  .ZN(_1673_)
);

NAND2_X1 _5858_ (
  .A1(_1672_),
  .A2(_1673_),
  .ZN(_1674_)
);

NAND2_X1 _5859_ (
  .A1(_4275_),
  .A2(_4278_),
  .ZN(_1675_)
);

NOR2_X1 _5860_ (
  .A1(_1636_),
  .A2(_1675_),
  .ZN(_1676_)
);

NAND2_X1 _5861_ (
  .A1(_1674_),
  .A2(_1676_),
  .ZN(_1677_)
);

INV_X1 _5862_ (
  .A(_1675_),
  .ZN(_1678_)
);

NAND2_X1 _5863_ (
  .A1(_1641_),
  .A2(_1678_),
  .ZN(_1679_)
);

INV_X1 _5864_ (
  .A(_4277_),
  .ZN(_1680_)
);

OAI21_X1 _5865_ (
  .A(_1680_),
  .B1(_1667_),
  .B2(_1659_),
  .ZN(_1681_)
);

INV_X1 _5866_ (
  .A(_1681_),
  .ZN(_1682_)
);

NAND2_X1 _5867_ (
  .A1(_1679_),
  .A2(_1682_),
  .ZN(_1683_)
);

INV_X1 _5868_ (
  .A(_1683_),
  .ZN(_1684_)
);

NAND4_X1 _5869_ (
  .A1(_1676_),
  .A2(_1613_),
  .A3(_1594_),
  .A4(_1570_),
  .ZN(_1685_)
);

NAND3_X1 _5870_ (
  .A1(_1677_),
  .A2(_1684_),
  .A3(_1685_),
  .ZN(_1686_)
);

NAND2_X1 _5871_ (
  .A1(_1686_),
  .A2(_4281_),
  .ZN(_1687_)
);

INV_X1 _5872_ (
  .A(_4281_),
  .ZN(_1688_)
);

NAND4_X1 _5873_ (
  .A1(_1677_),
  .A2(_1685_),
  .A3(_1684_),
  .A4(_1688_),
  .ZN(_1689_)
);

NAND3_X1 _5874_ (
  .A1(_1687_),
  .A2(_1689_),
  .A3(_1669_),
  .ZN(_1690_)
);

NAND2_X1 _5875_ (
  .A1(_1490_),
  .A2(\s_pipe[1][22] ),
  .ZN(_1691_)
);

NAND2_X1 _5876_ (
  .A1(_1690_),
  .A2(_1691_),
  .ZN(_0202_)
);

NAND2_X1 _5877_ (
  .A1(_4278_),
  .A2(_4281_),
  .ZN(_1692_)
);

OR2_X2 _5878_ (
  .A1(_1692_),
  .A2(_1654_),
  .ZN(_1693_)
);

INV_X1 _5879_ (
  .A(_1693_),
  .ZN(_1694_)
);

NAND2_X1 _5880_ (
  .A1(_1627_),
  .A2(_1694_),
  .ZN(_1695_)
);

INV_X1 _5881_ (
  .A(_4280_),
  .ZN(_1696_)
);

OAI21_X1 _5882_ (
  .A(_1696_),
  .B1(_1688_),
  .B2(_1680_),
  .ZN(_1697_)
);

INV_X1 _5883_ (
  .A(_1697_),
  .ZN(_1698_)
);

OAI21_X1 _5884_ (
  .A(_1698_),
  .B1(_1661_),
  .B2(_1692_),
  .ZN(_1699_)
);

INV_X1 _5885_ (
  .A(_1699_),
  .ZN(_1700_)
);

INV_X1 _5886_ (
  .A(_4284_),
  .ZN(_1701_)
);

NAND2_X1 _5887_ (
  .A1(_1603_),
  .A2(_1621_),
  .ZN(_1702_)
);

NOR2_X1 _5888_ (
  .A1(_1693_),
  .A2(_1702_),
  .ZN(_1703_)
);

NAND2_X1 _5889_ (
  .A1(_1584_),
  .A2(_1703_),
  .ZN(_1704_)
);

NAND4_X1 _5890_ (
  .A1(_1695_),
  .A2(_1700_),
  .A3(_1701_),
  .A4(_1704_),
  .ZN(_1705_)
);

NAND3_X1 _5891_ (
  .A1(_1695_),
  .A2(_1700_),
  .A3(_1704_),
  .ZN(_1706_)
);

NAND2_X1 _5892_ (
  .A1(_1706_),
  .A2(_4284_),
  .ZN(_1707_)
);

NAND3_X1 _5893_ (
  .A1(_1705_),
  .A2(_1707_),
  .A3(_1669_),
  .ZN(_1708_)
);

BUF_X4 _5894_ (
  .A(_1337_),
  .Z(_1709_)
);

NAND2_X1 _5895_ (
  .A1(_1709_),
  .A2(\s_pipe[1][23] ),
  .ZN(_1710_)
);

NAND2_X1 _5896_ (
  .A1(_1708_),
  .A2(_1710_),
  .ZN(_0203_)
);

NAND2_X1 _5897_ (
  .A1(_4281_),
  .A2(_4284_),
  .ZN(_1711_)
);

OR2_X2 _5898_ (
  .A1(_1711_),
  .A2(_1675_),
  .ZN(_1712_)
);

INV_X1 _5899_ (
  .A(_1712_),
  .ZN(_1713_)
);

NAND2_X1 _5900_ (
  .A1(_1643_),
  .A2(_1713_),
  .ZN(_1714_)
);

INV_X1 _5901_ (
  .A(_4283_),
  .ZN(_1715_)
);

OAI21_X1 _5902_ (
  .A(_1715_),
  .B1(_1701_),
  .B2(_1696_),
  .ZN(_1716_)
);

INV_X1 _5903_ (
  .A(_1716_),
  .ZN(_1717_)
);

OAI21_X1 _5904_ (
  .A(_1717_),
  .B1(_1682_),
  .B2(_1711_),
  .ZN(_1718_)
);

INV_X1 _5905_ (
  .A(_1718_),
  .ZN(_1719_)
);

NAND2_X1 _5906_ (
  .A1(_1613_),
  .A2(_1637_),
  .ZN(_1720_)
);

NOR2_X1 _5907_ (
  .A1(_1712_),
  .A2(_1720_),
  .ZN(_1721_)
);

NAND2_X1 _5908_ (
  .A1(_1596_),
  .A2(_1721_),
  .ZN(_1722_)
);

NAND4_X1 _5909_ (
  .A1(_1714_),
  .A2(_1719_),
  .A3(z[23]),
  .A4(_1722_),
  .ZN(_1723_)
);

NAND3_X1 _5910_ (
  .A1(_1714_),
  .A2(_1719_),
  .A3(_1722_),
  .ZN(_1724_)
);

INV_X1 _5911_ (
  .A(z[23]),
  .ZN(_1725_)
);

NAND2_X1 _5912_ (
  .A1(_1724_),
  .A2(_1725_),
  .ZN(_1726_)
);

NAND3_X1 _5913_ (
  .A1(_1723_),
  .A2(_1726_),
  .A3(_1669_),
  .ZN(_1727_)
);

BUF_X2 _5914_ (
  .A(_1340_),
  .Z(_1728_)
);

NAND2_X1 _5915_ (
  .A1(_1728_),
  .A2(\s_pipe[1][24] ),
  .ZN(_1729_)
);

NAND2_X1 _5916_ (
  .A1(_1727_),
  .A2(_1729_),
  .ZN(_0204_)
);

BUF_X2 _6049_ (
  .A(_1340_),
  .Z(_1859_)
);

MUX2_X1 _6052_ (
  .A(\q_pipe[1] ),
  .B(_0111_),
  .S(_1336_),
  .Z(_0209_)
);

BUF_X2 _6053_ (
  .A(_1335_),
  .Z(_1861_)
);

MUX2_X1 _6054_ (
  .A(q[0]),
  .B(_0122_),
  .S(_1861_),
  .Z(_0210_)
);

NAND2_X1 _6055_ (
  .A1(_1338_),
  .A2(q[1]),
  .ZN(_1862_)
);

INV_X1 _6056_ (
  .A(\q_pipe[11][0] ),
  .ZN(_1863_)
);

OAI21_X1 _6057_ (
  .A(_1862_),
  .B1(_1524_),
  .B2(_1863_),
  .ZN(_0211_)
);

NAND2_X1 _6058_ (
  .A1(_1338_),
  .A2(q[2]),
  .ZN(_1864_)
);

BUF_X2 _6059_ (
  .A(_1522_),
  .Z(_1865_)
);

INV_X1 _6060_ (
  .A(\q_pipe[11][1] ),
  .ZN(_1866_)
);

OAI21_X1 _6061_ (
  .A(_1864_),
  .B1(_1865_),
  .B2(_1866_),
  .ZN(_0212_)
);

NAND2_X1 _6062_ (
  .A1(_1338_),
  .A2(q[3]),
  .ZN(_1867_)
);

INV_X1 _6063_ (
  .A(\q_pipe[11][2] ),
  .ZN(_1868_)
);

OAI21_X1 _6064_ (
  .A(_1867_),
  .B1(_1865_),
  .B2(_1868_),
  .ZN(_0213_)
);

NAND2_X1 _6065_ (
  .A1(_1338_),
  .A2(q[4]),
  .ZN(_1869_)
);

INV_X1 _6066_ (
  .A(\q_pipe[11][3] ),
  .ZN(_1870_)
);

OAI21_X1 _6067_ (
  .A(_1869_),
  .B1(_1865_),
  .B2(_1870_),
  .ZN(_0214_)
);

NAND2_X1 _6068_ (
  .A1(_1338_),
  .A2(q[5]),
  .ZN(_1871_)
);

INV_X1 _6069_ (
  .A(\q_pipe[11][4] ),
  .ZN(_1872_)
);

OAI21_X1 _6070_ (
  .A(_1871_),
  .B1(_1865_),
  .B2(_1872_),
  .ZN(_0215_)
);

NAND2_X1 _6071_ (
  .A1(_1522_),
  .A2(q[6]),
  .ZN(_1873_)
);

INV_X1 _6072_ (
  .A(\q_pipe[11][5] ),
  .ZN(_1874_)
);

OAI21_X1 _6073_ (
  .A(_1873_),
  .B1(_1865_),
  .B2(_1874_),
  .ZN(_0216_)
);

NAND2_X1 _6074_ (
  .A1(_1338_),
  .A2(q[7]),
  .ZN(_1875_)
);

INV_X1 _6075_ (
  .A(\q_pipe[11][6] ),
  .ZN(_1876_)
);

OAI21_X1 _6076_ (
  .A(_1875_),
  .B1(_1524_),
  .B2(_1876_),
  .ZN(_0217_)
);

NAND2_X1 _6077_ (
  .A1(_1338_),
  .A2(q[8]),
  .ZN(_1877_)
);

INV_X1 _6078_ (
  .A(\q_pipe[11][7] ),
  .ZN(_1878_)
);

OAI21_X1 _6079_ (
  .A(_1877_),
  .B1(_1865_),
  .B2(_1878_),
  .ZN(_0218_)
);

NAND2_X1 _6080_ (
  .A1(_1338_),
  .A2(q[9]),
  .ZN(_1879_)
);

INV_X1 _6081_ (
  .A(\q_pipe[11][8] ),
  .ZN(_1880_)
);

OAI21_X1 _6082_ (
  .A(_1879_),
  .B1(_1524_),
  .B2(_1880_),
  .ZN(_0219_)
);

BUF_X1 _6083_ (
  .A(_1337_),
  .Z(_1881_)
);

NAND2_X1 _6084_ (
  .A1(_1881_),
  .A2(q[10]),
  .ZN(_1882_)
);

INV_X1 _6085_ (
  .A(\q_pipe[11][9] ),
  .ZN(_1883_)
);

OAI21_X1 _6086_ (
  .A(_1882_),
  .B1(_1524_),
  .B2(_1883_),
  .ZN(_0220_)
);

NAND2_X1 _6087_ (
  .A1(_1881_),
  .A2(q[11]),
  .ZN(_1884_)
);

INV_X1 _6088_ (
  .A(\q_pipe[11][10] ),
  .ZN(_1885_)
);

OAI21_X1 _6089_ (
  .A(_1884_),
  .B1(_1524_),
  .B2(_1885_),
  .ZN(_0221_)
);

NOR2_X1 _6099_ (
  .A1(_1337_),
  .A2(d[0]),
  .ZN(_1893_)
);

BUF_X2 _6105_ (
  .A(_1335_),
  .Z(_1897_)
);

BUF_X2 _6108_ (
  .A(_1335_),
  .Z(_1898_)
);

BUF_X2 _6116_ (
  .A(_1446_),
  .Z(_1899_)
);

BUF_X2 _6118_ (
  .A(_1350_),
  .Z(_1901_)
);

BUF_X2 _6154_ (
  .A(_1335_),
  .Z(_1933_)
);

BUF_X2 _6157_ (
  .A(_1335_),
  .Z(_1934_)
);

INV_X1 _6166_ (
  .A(\d_pipe[1][12] ),
  .ZN(_1936_)
);

AOI21_X1 _6167_ (
  .A(_1893_),
  .B1(_1936_),
  .B2(_1865_),
  .ZN(_0248_)
);

BUF_X2 _6168_ (
  .A(_1526_),
  .Z(_1937_)
);

NAND2_X1 _6169_ (
  .A1(d[1]),
  .A2(_1937_),
  .ZN(_1938_)
);

OAI21_X1 _6170_ (
  .A(_1938_),
  .B1(_0672_),
  .B2(_1535_),
  .ZN(_0249_)
);

NAND2_X1 _6171_ (
  .A1(d[2]),
  .A2(_1937_),
  .ZN(_1939_)
);

OAI21_X1 _6172_ (
  .A(_1939_),
  .B1(_0671_),
  .B2(_1535_),
  .ZN(_0250_)
);

NAND2_X1 _6173_ (
  .A1(d[3]),
  .A2(_1937_),
  .ZN(_1940_)
);

OAI21_X1 _6174_ (
  .A(_1940_),
  .B1(_0675_),
  .B2(_1535_),
  .ZN(_0251_)
);

NAND2_X1 _6175_ (
  .A1(d[4]),
  .A2(_1937_),
  .ZN(_1941_)
);

OAI21_X1 _6176_ (
  .A(_1941_),
  .B1(_0810_),
  .B2(_1535_),
  .ZN(_0252_)
);

BUF_X2 _6177_ (
  .A(_1526_),
  .Z(_1942_)
);

NAND2_X1 _6178_ (
  .A1(d[5]),
  .A2(_1942_),
  .ZN(_1943_)
);

BUF_X2 _6179_ (
  .A(_1426_),
  .Z(_1944_)
);

OAI21_X1 _6180_ (
  .A(_1943_),
  .B1(_0812_),
  .B2(_1944_),
  .ZN(_0253_)
);

NAND2_X1 _6181_ (
  .A1(d[6]),
  .A2(_1942_),
  .ZN(_1945_)
);

OAI21_X1 _6182_ (
  .A(_1945_),
  .B1(_0817_),
  .B2(_1944_),
  .ZN(_0254_)
);

NAND2_X1 _6183_ (
  .A1(d[7]),
  .A2(_1942_),
  .ZN(_1946_)
);

OAI21_X1 _6184_ (
  .A(_1946_),
  .B1(_0823_),
  .B2(_1944_),
  .ZN(_0255_)
);

NAND2_X1 _6185_ (
  .A1(d[8]),
  .A2(_1942_),
  .ZN(_1947_)
);

OAI21_X1 _6186_ (
  .A(_1947_),
  .B1(_0830_),
  .B2(_1944_),
  .ZN(_0256_)
);

NAND2_X1 _6187_ (
  .A1(d[9]),
  .A2(_1942_),
  .ZN(_1948_)
);

OAI21_X1 _6188_ (
  .A(_1948_),
  .B1(_0838_),
  .B2(_1944_),
  .ZN(_0257_)
);

BUF_X2 _6189_ (
  .A(_1526_),
  .Z(_1949_)
);

NAND2_X1 _6190_ (
  .A1(d[10]),
  .A2(_1949_),
  .ZN(_1950_)
);

OAI21_X1 _6191_ (
  .A(_1950_),
  .B1(_0843_),
  .B2(_1533_),
  .ZN(_0258_)
);

NAND2_X1 _6192_ (
  .A1(d[11]),
  .A2(_1949_),
  .ZN(_1951_)
);

OAI21_X1 _6193_ (
  .A(_1951_),
  .B1(_0851_),
  .B2(_1533_),
  .ZN(_0259_)
);

BUF_X2 _6194_ (
  .A(_1346_),
  .Z(_1952_)
);

MUX2_X1 _6195_ (
  .A(\d_pipe[4][12] ),
  .B(\d_pipe[3][12] ),
  .S(_1952_),
  .Z(_0260_)
);

NAND2_X1 _6196_ (
  .A1(\d_pipe[3][13] ),
  .A2(_1949_),
  .ZN(_1953_)
);

OAI21_X1 _6197_ (
  .A(_1953_),
  .B1(_1275_),
  .B2(_1533_),
  .ZN(_0261_)
);

NAND2_X1 _6198_ (
  .A1(\d_pipe[3][14] ),
  .A2(_1949_),
  .ZN(_1954_)
);

OAI21_X1 _6199_ (
  .A(_1954_),
  .B1(_1274_),
  .B2(_1533_),
  .ZN(_0262_)
);

NAND2_X1 _6200_ (
  .A1(\d_pipe[3][15] ),
  .A2(_1949_),
  .ZN(_1955_)
);

OAI21_X1 _6201_ (
  .A(_1955_),
  .B1(_1278_),
  .B2(_1533_),
  .ZN(_0263_)
);

BUF_X2 _6202_ (
  .A(_1446_),
  .Z(_1956_)
);

NAND2_X1 _6203_ (
  .A1(_0756_),
  .A2(_1956_),
  .ZN(_1957_)
);

BUF_X2 _6204_ (
  .A(_1426_),
  .Z(_1958_)
);

OAI21_X1 _6205_ (
  .A(_1957_),
  .B1(_1298_),
  .B2(_1958_),
  .ZN(_0264_)
);

NAND2_X1 _6206_ (
  .A1(_0763_),
  .A2(_1956_),
  .ZN(_1959_)
);

OAI21_X1 _6207_ (
  .A(_1959_),
  .B1(_1288_),
  .B2(_1958_),
  .ZN(_0265_)
);

NAND2_X1 _6208_ (
  .A1(\d_pipe[3][18] ),
  .A2(_1956_),
  .ZN(_1960_)
);

OAI21_X1 _6209_ (
  .A(_1960_),
  .B1(_1294_),
  .B2(_1958_),
  .ZN(_0266_)
);

NAND2_X1 _6210_ (
  .A1(\d_pipe[3][19] ),
  .A2(_1956_),
  .ZN(_1961_)
);

OAI21_X1 _6211_ (
  .A(_1961_),
  .B1(_1301_),
  .B2(_1958_),
  .ZN(_0267_)
);

BUF_X2 _6212_ (
  .A(_1526_),
  .Z(_1962_)
);

NAND2_X1 _6213_ (
  .A1(\d_pipe[3][20] ),
  .A2(_1962_),
  .ZN(_1963_)
);

OAI21_X1 _6214_ (
  .A(_1963_),
  .B1(_1308_),
  .B2(_1958_),
  .ZN(_0268_)
);

NAND2_X1 _6215_ (
  .A1(\d_pipe[3][21] ),
  .A2(_1937_),
  .ZN(_1964_)
);

OAI21_X1 _6216_ (
  .A(_1964_),
  .B1(_1326_),
  .B2(_1531_),
  .ZN(_0269_)
);

NAND2_X1 _6217_ (
  .A1(\d_pipe[3][22] ),
  .A2(_1937_),
  .ZN(_1965_)
);

OAI21_X1 _6218_ (
  .A(_1965_),
  .B1(_1322_),
  .B2(_1531_),
  .ZN(_0270_)
);

BUF_X2 _6219_ (
  .A(_1526_),
  .Z(_1966_)
);

NAND2_X1 _6220_ (
  .A1(\d_pipe[3][23] ),
  .A2(_1966_),
  .ZN(_1967_)
);

OAI21_X1 _6221_ (
  .A(_1967_),
  .B1(_1331_),
  .B2(_1531_),
  .ZN(_0271_)
);

MUX2_X1 _6222_ (
  .A(\d_pipe[5][12] ),
  .B(\d_pipe[4][12] ),
  .S(_1952_),
  .Z(_0272_)
);

NAND2_X1 _6223_ (
  .A1(\d_pipe[4][13] ),
  .A2(_1966_),
  .ZN(_1968_)
);

OAI21_X1 _6224_ (
  .A(_1968_),
  .B1(_1212_),
  .B2(_1531_),
  .ZN(_0273_)
);

NAND2_X1 _6225_ (
  .A1(\d_pipe[4][14] ),
  .A2(_1966_),
  .ZN(_1969_)
);

BUF_X2 _6226_ (
  .A(_1426_),
  .Z(_1970_)
);

OAI21_X1 _6227_ (
  .A(_1969_),
  .B1(_1211_),
  .B2(_1970_),
  .ZN(_0274_)
);

NAND2_X1 _6228_ (
  .A1(\d_pipe[4][15] ),
  .A2(_1966_),
  .ZN(_1971_)
);

OAI21_X1 _6229_ (
  .A(_1971_),
  .B1(_1215_),
  .B2(_1970_),
  .ZN(_0275_)
);

NAND2_X1 _6230_ (
  .A1(_1283_),
  .A2(_1966_),
  .ZN(_1972_)
);

OAI21_X1 _6231_ (
  .A(_1972_),
  .B1(_1235_),
  .B2(_1970_),
  .ZN(_0276_)
);

NAND2_X1 _6232_ (
  .A1(_1287_),
  .A2(_1962_),
  .ZN(_1973_)
);

OAI21_X1 _6233_ (
  .A(_1973_),
  .B1(_1225_),
  .B2(_1970_),
  .ZN(_0277_)
);

NAND2_X1 _6234_ (
  .A1(\d_pipe[4][18] ),
  .A2(_1962_),
  .ZN(_1974_)
);

OAI21_X1 _6235_ (
  .A(_1974_),
  .B1(_1231_),
  .B2(_1970_),
  .ZN(_0278_)
);

NAND2_X1 _6236_ (
  .A1(\d_pipe[4][19] ),
  .A2(_1962_),
  .ZN(_1975_)
);

OAI21_X1 _6237_ (
  .A(_1975_),
  .B1(_1238_),
  .B2(_1529_),
  .ZN(_0279_)
);

BUF_X2 _6238_ (
  .A(_1347_),
  .Z(_1976_)
);

NAND2_X1 _6239_ (
  .A1(\d_pipe[4][20] ),
  .A2(_1976_),
  .ZN(_1977_)
);

OAI21_X1 _6240_ (
  .A(_1977_),
  .B1(_1245_),
  .B2(_1529_),
  .ZN(_0280_)
);

NAND2_X1 _6241_ (
  .A1(_1314_),
  .A2(_1962_),
  .ZN(_1978_)
);

OAI21_X1 _6242_ (
  .A(_1978_),
  .B1(_1263_),
  .B2(_1529_),
  .ZN(_0281_)
);

BUF_X2 _6243_ (
  .A(_1526_),
  .Z(_1979_)
);

NAND2_X1 _6244_ (
  .A1(\d_pipe[4][22] ),
  .A2(_1979_),
  .ZN(_1980_)
);

OAI21_X1 _6245_ (
  .A(_1980_),
  .B1(_1259_),
  .B2(_1529_),
  .ZN(_0282_)
);

NAND2_X1 _6246_ (
  .A1(\d_pipe[4][23] ),
  .A2(_1979_),
  .ZN(_1981_)
);

OAI21_X1 _6247_ (
  .A(_1981_),
  .B1(_1268_),
  .B2(_1529_),
  .ZN(_0283_)
);

MUX2_X1 _6248_ (
  .A(\d_pipe[6][12] ),
  .B(\d_pipe[5][12] ),
  .S(_1934_),
  .Z(_0284_)
);

NAND2_X1 _6249_ (
  .A1(\d_pipe[5][13] ),
  .A2(_1979_),
  .ZN(_1982_)
);

OAI21_X1 _6250_ (
  .A(_1982_),
  .B1(_1152_),
  .B2(_1427_),
  .ZN(_0285_)
);

NAND2_X1 _6251_ (
  .A1(\d_pipe[5][14] ),
  .A2(_1979_),
  .ZN(_1983_)
);

OAI21_X1 _6252_ (
  .A(_1983_),
  .B1(_1151_),
  .B2(_1427_),
  .ZN(_0286_)
);

NAND2_X1 _6253_ (
  .A1(\d_pipe[5][15] ),
  .A2(_1979_),
  .ZN(_1984_)
);

OAI21_X1 _6254_ (
  .A(_1984_),
  .B1(_1155_),
  .B2(_1427_),
  .ZN(_0287_)
);

NAND2_X1 _6255_ (
  .A1(_1220_),
  .A2(_1558_),
  .ZN(_1985_)
);

OAI21_X1 _6256_ (
  .A(_1985_),
  .B1(_1164_),
  .B2(_1427_),
  .ZN(_0288_)
);

NAND2_X1 _6257_ (
  .A1(_1224_),
  .A2(_1558_),
  .ZN(_1986_)
);

OAI21_X1 _6258_ (
  .A(_1986_),
  .B1(_1166_),
  .B2(_1427_),
  .ZN(_0289_)
);

NAND2_X1 _6259_ (
  .A1(\d_pipe[5][18] ),
  .A2(_1976_),
  .ZN(_1987_)
);

BUF_X2 _6260_ (
  .A(_1446_),
  .Z(_1988_)
);

OAI21_X1 _6261_ (
  .A(_1987_),
  .B1(_1171_),
  .B2(_1988_),
  .ZN(_0290_)
);

NAND2_X1 _6262_ (
  .A1(\d_pipe[5][19] ),
  .A2(_1558_),
  .ZN(_1989_)
);

OAI21_X1 _6263_ (
  .A(_1989_),
  .B1(_1177_),
  .B2(_1988_),
  .ZN(_0291_)
);

NAND2_X1 _6264_ (
  .A1(\d_pipe[5][20] ),
  .A2(_1558_),
  .ZN(_1990_)
);

OAI21_X1 _6265_ (
  .A(_1990_),
  .B1(_1184_),
  .B2(_1988_),
  .ZN(_0292_)
);

NAND2_X1 _6266_ (
  .A1(_1251_),
  .A2(_1537_),
  .ZN(_1991_)
);

OAI21_X1 _6267_ (
  .A(_1991_),
  .B1(_1192_),
  .B2(_1988_),
  .ZN(_0293_)
);

NAND2_X1 _6268_ (
  .A1(\d_pipe[5][22] ),
  .A2(_1537_),
  .ZN(_1992_)
);

OAI21_X1 _6269_ (
  .A(_1992_),
  .B1(_1197_),
  .B2(_1988_),
  .ZN(_0294_)
);

NAND2_X1 _6270_ (
  .A1(\d_pipe[5][23] ),
  .A2(_1537_),
  .ZN(_1993_)
);

BUF_X2 _6271_ (
  .A(_1446_),
  .Z(_1994_)
);

OAI21_X1 _6272_ (
  .A(_1993_),
  .B1(_1205_),
  .B2(_1994_),
  .ZN(_0295_)
);

MUX2_X1 _6273_ (
  .A(\d_pipe[7][12] ),
  .B(\d_pipe[6][12] ),
  .S(_1934_),
  .Z(_0296_)
);

NAND2_X1 _6274_ (
  .A1(\d_pipe[6][13] ),
  .A2(_1527_),
  .ZN(_1995_)
);

OAI21_X1 _6275_ (
  .A(_1995_),
  .B1(_1091_),
  .B2(_1994_),
  .ZN(_0297_)
);

NAND2_X1 _6276_ (
  .A1(\d_pipe[6][14] ),
  .A2(_1527_),
  .ZN(_1996_)
);

OAI21_X1 _6277_ (
  .A(_1996_),
  .B1(_1090_),
  .B2(_1994_),
  .ZN(_0298_)
);

NAND2_X1 _6278_ (
  .A1(\d_pipe[6][15] ),
  .A2(_1976_),
  .ZN(_1997_)
);

OAI21_X1 _6279_ (
  .A(_1997_),
  .B1(_1094_),
  .B2(_1994_),
  .ZN(_0299_)
);

NAND2_X1 _6280_ (
  .A1(_1160_),
  .A2(_1976_),
  .ZN(_1998_)
);

OAI21_X1 _6281_ (
  .A(_1998_),
  .B1(_1103_),
  .B2(_1546_),
  .ZN(_0300_)
);

NAND2_X1 _6282_ (
  .A1(_1165_),
  .A2(_1976_),
  .ZN(_1999_)
);

OAI21_X1 _6283_ (
  .A(_1999_),
  .B1(_1107_),
  .B2(_1994_),
  .ZN(_0301_)
);

NAND2_X1 _6284_ (
  .A1(\d_pipe[6][18] ),
  .A2(_1558_),
  .ZN(_2000_)
);

OAI21_X1 _6285_ (
  .A(_2000_),
  .B1(_1111_),
  .B2(_1546_),
  .ZN(_0302_)
);

BUF_X2 _6286_ (
  .A(_1446_),
  .Z(_2001_)
);

NAND2_X1 _6287_ (
  .A1(\d_pipe[6][19] ),
  .A2(_2001_),
  .ZN(_2002_)
);

OAI21_X1 _6288_ (
  .A(_2002_),
  .B1(_1127_),
  .B2(_1552_),
  .ZN(_0303_)
);

NAND2_X1 _6289_ (
  .A1(\d_pipe[6][20] ),
  .A2(_1976_),
  .ZN(_2003_)
);

OAI21_X1 _6290_ (
  .A(_2003_),
  .B1(_1123_),
  .B2(_1994_),
  .ZN(_0304_)
);

NAND2_X1 _6291_ (
  .A1(\d_pipe[6][21] ),
  .A2(_1976_),
  .ZN(_2004_)
);

OAI21_X1 _6292_ (
  .A(_2004_),
  .B1(_1132_),
  .B2(_1994_),
  .ZN(_0305_)
);

NAND2_X1 _6293_ (
  .A1(\d_pipe[6][22] ),
  .A2(_1527_),
  .ZN(_2005_)
);

OAI21_X1 _6294_ (
  .A(_2005_),
  .B1(_1137_),
  .B2(_1994_),
  .ZN(_0306_)
);

NAND2_X1 _6295_ (
  .A1(\d_pipe[6][23] ),
  .A2(_1527_),
  .ZN(_2006_)
);

OAI21_X1 _6296_ (
  .A(_2006_),
  .B1(_1145_),
  .B2(_1994_),
  .ZN(_0307_)
);

BUF_X2 _6297_ (
  .A(_1346_),
  .Z(_2007_)
);

MUX2_X1 _6298_ (
  .A(\d_pipe[8][12] ),
  .B(\d_pipe[7][12] ),
  .S(_2007_),
  .Z(_0308_)
);

NAND2_X1 _6299_ (
  .A1(\d_pipe[7][13] ),
  .A2(_1527_),
  .ZN(_2008_)
);

OAI21_X1 _6300_ (
  .A(_2008_),
  .B1(_1030_),
  .B2(_1994_),
  .ZN(_0309_)
);

NAND2_X1 _6301_ (
  .A1(\d_pipe[7][14] ),
  .A2(_1537_),
  .ZN(_2009_)
);

OAI21_X1 _6302_ (
  .A(_2009_),
  .B1(_1029_),
  .B2(_1988_),
  .ZN(_0310_)
);

NAND2_X1 _6303_ (
  .A1(\d_pipe[7][15] ),
  .A2(_1537_),
  .ZN(_2010_)
);

OAI21_X1 _6304_ (
  .A(_2010_),
  .B1(_1033_),
  .B2(_1988_),
  .ZN(_0311_)
);

NAND2_X1 _6305_ (
  .A1(_1099_),
  .A2(_1544_),
  .ZN(_2011_)
);

OAI21_X1 _6306_ (
  .A(_2011_),
  .B1(_1042_),
  .B2(_1988_),
  .ZN(_0312_)
);

NAND2_X1 _6307_ (
  .A1(_1106_),
  .A2(_1976_),
  .ZN(_2012_)
);

OAI21_X1 _6308_ (
  .A(_2012_),
  .B1(_1046_),
  .B2(_1988_),
  .ZN(_0313_)
);

NAND2_X1 _6309_ (
  .A1(\d_pipe[7][18] ),
  .A2(_1976_),
  .ZN(_2013_)
);

OAI21_X1 _6310_ (
  .A(_2013_),
  .B1(_1050_),
  .B2(_1988_),
  .ZN(_0314_)
);

NAND2_X1 _6311_ (
  .A1(\d_pipe[7][19] ),
  .A2(_1558_),
  .ZN(_2014_)
);

OAI21_X1 _6312_ (
  .A(_2014_),
  .B1(_1066_),
  .B2(_1427_),
  .ZN(_0315_)
);

NAND2_X1 _6313_ (
  .A1(\d_pipe[7][20] ),
  .A2(_1558_),
  .ZN(_2015_)
);

OAI21_X1 _6314_ (
  .A(_2015_),
  .B1(_1062_),
  .B2(_1427_),
  .ZN(_0316_)
);

NAND2_X1 _6315_ (
  .A1(\d_pipe[7][21] ),
  .A2(_1558_),
  .ZN(_2016_)
);

OAI21_X1 _6316_ (
  .A(_2016_),
  .B1(_1071_),
  .B2(_1427_),
  .ZN(_0317_)
);

NAND2_X1 _6317_ (
  .A1(\d_pipe[7][22] ),
  .A2(_1979_),
  .ZN(_2017_)
);

OAI21_X1 _6318_ (
  .A(_2017_),
  .B1(_1076_),
  .B2(_1546_),
  .ZN(_0318_)
);

NAND2_X1 _6319_ (
  .A1(\d_pipe[7][23] ),
  .A2(_1979_),
  .ZN(_2018_)
);

OAI21_X1 _6320_ (
  .A(_2018_),
  .B1(_1084_),
  .B2(_1427_),
  .ZN(_0319_)
);

MUX2_X1 _6321_ (
  .A(\d_pipe[9][12] ),
  .B(\d_pipe[8][12] ),
  .S(_1934_),
  .Z(_0320_)
);

NAND2_X1 _6322_ (
  .A1(\d_pipe[8][13] ),
  .A2(_1979_),
  .ZN(_2019_)
);

OAI21_X1 _6323_ (
  .A(_2019_),
  .B1(_0976_),
  .B2(_1529_),
  .ZN(_0321_)
);

NAND2_X1 _6324_ (
  .A1(\d_pipe[8][14] ),
  .A2(_1979_),
  .ZN(_2020_)
);

OAI21_X1 _6325_ (
  .A(_2020_),
  .B1(_0679_),
  .B2(_1529_),
  .ZN(_0322_)
);

NAND2_X1 _6326_ (
  .A1(\d_pipe[8][15] ),
  .A2(_1979_),
  .ZN(_2021_)
);

OAI21_X1 _6327_ (
  .A(_2021_),
  .B1(_0680_),
  .B2(_1529_),
  .ZN(_0323_)
);

NAND2_X1 _6328_ (
  .A1(_1038_),
  .A2(_1962_),
  .ZN(_2022_)
);

OAI21_X1 _6329_ (
  .A(_2022_),
  .B1(_0982_),
  .B2(_1529_),
  .ZN(_0324_)
);

NAND2_X1 _6330_ (
  .A1(_1045_),
  .A2(_1962_),
  .ZN(_2023_)
);

OAI21_X1 _6331_ (
  .A(_2023_),
  .B1(_0984_),
  .B2(_1970_),
  .ZN(_0325_)
);

NAND2_X1 _6332_ (
  .A1(\d_pipe[8][18] ),
  .A2(_1962_),
  .ZN(_2024_)
);

OAI21_X1 _6333_ (
  .A(_2024_),
  .B1(_0989_),
  .B2(_1970_),
  .ZN(_0326_)
);

NAND2_X1 _6334_ (
  .A1(\d_pipe[8][19] ),
  .A2(_1962_),
  .ZN(_2025_)
);

OAI21_X1 _6335_ (
  .A(_2025_),
  .B1(_0995_),
  .B2(_1970_),
  .ZN(_0327_)
);

NAND2_X1 _6336_ (
  .A1(\d_pipe[8][20] ),
  .A2(_1962_),
  .ZN(_2026_)
);

OAI21_X1 _6337_ (
  .A(_2026_),
  .B1(_1002_),
  .B2(_1970_),
  .ZN(_0328_)
);

NAND2_X1 _6338_ (
  .A1(\d_pipe[8][21] ),
  .A2(_1966_),
  .ZN(_2027_)
);

OAI21_X1 _6339_ (
  .A(_2027_),
  .B1(_1010_),
  .B2(_1970_),
  .ZN(_0329_)
);

NAND2_X1 _6340_ (
  .A1(\d_pipe[8][22] ),
  .A2(_1966_),
  .ZN(_2028_)
);

OAI21_X1 _6341_ (
  .A(_2028_),
  .B1(_1015_),
  .B2(_1531_),
  .ZN(_0330_)
);

NAND2_X1 _6342_ (
  .A1(\d_pipe[8][23] ),
  .A2(_1966_),
  .ZN(_2029_)
);

OAI21_X1 _6343_ (
  .A(_2029_),
  .B1(_1023_),
  .B2(_1531_),
  .ZN(_0331_)
);

MUX2_X1 _6344_ (
  .A(\d_pipe[10][12] ),
  .B(\d_pipe[9][12] ),
  .S(_1934_),
  .Z(_0332_)
);

NAND2_X1 _6345_ (
  .A1(_3714_),
  .A2(_1966_),
  .ZN(_2030_)
);

OAI21_X1 _6346_ (
  .A(_2030_),
  .B1(_0918_),
  .B2(_1531_),
  .ZN(_0333_)
);

NAND2_X1 _6347_ (
  .A1(_3715_),
  .A2(_1966_),
  .ZN(_2031_)
);

OAI21_X1 _6348_ (
  .A(_2031_),
  .B1(_0917_),
  .B2(_1546_),
  .ZN(_0334_)
);

NAND2_X1 _6349_ (
  .A1(_3716_),
  .A2(_1937_),
  .ZN(_2032_)
);

OAI21_X1 _6350_ (
  .A(_2032_),
  .B1(_0921_),
  .B2(_1531_),
  .ZN(_0335_)
);

NAND2_X1 _6351_ (
  .A1(_0682_),
  .A2(_1956_),
  .ZN(_2033_)
);

OAI21_X1 _6352_ (
  .A(_2033_),
  .B1(_0930_),
  .B2(_1958_),
  .ZN(_0336_)
);

NAND2_X1 _6353_ (
  .A1(_0983_),
  .A2(_1956_),
  .ZN(_2034_)
);

OAI21_X1 _6354_ (
  .A(_2034_),
  .B1(_0932_),
  .B2(_1958_),
  .ZN(_0337_)
);

NAND2_X1 _6355_ (
  .A1(_3719_),
  .A2(_1956_),
  .ZN(_2035_)
);

OAI21_X1 _6356_ (
  .A(_2035_),
  .B1(_0937_),
  .B2(_1958_),
  .ZN(_0338_)
);

NAND2_X1 _6357_ (
  .A1(_3720_),
  .A2(_1956_),
  .ZN(_2036_)
);

OAI21_X1 _6358_ (
  .A(_2036_),
  .B1(_0943_),
  .B2(_1958_),
  .ZN(_0339_)
);

NAND2_X1 _6359_ (
  .A1(_3721_),
  .A2(_1956_),
  .ZN(_2037_)
);

OAI21_X1 _6360_ (
  .A(_2037_),
  .B1(_0950_),
  .B2(_1958_),
  .ZN(_0340_)
);

NAND2_X1 _6361_ (
  .A1(_3722_),
  .A2(_1956_),
  .ZN(_2038_)
);

OAI21_X1 _6362_ (
  .A(_2038_),
  .B1(_0958_),
  .B2(_1533_),
  .ZN(_0341_)
);

NAND2_X1 _6363_ (
  .A1(_3712_),
  .A2(_1949_),
  .ZN(_2039_)
);

OAI21_X1 _6364_ (
  .A(_2039_),
  .B1(_0963_),
  .B2(_1533_),
  .ZN(_0342_)
);

NAND2_X1 _6365_ (
  .A1(_3713_),
  .A2(_1949_),
  .ZN(_2040_)
);

OAI21_X1 _6366_ (
  .A(_2040_),
  .B1(_0971_),
  .B2(_1533_),
  .ZN(_0343_)
);

BUF_X4 _6367_ (
  .A(_1347_),
  .Z(_2041_)
);

MUX2_X1 _6368_ (
  .A(\d_pipe[11][12] ),
  .B(\d_pipe[10][12] ),
  .S(_2041_),
  .Z(_0344_)
);

NAND2_X1 _6369_ (
  .A1(\d_pipe[10][13] ),
  .A2(_1949_),
  .ZN(_2042_)
);

OAI21_X1 _6370_ (
  .A(_2042_),
  .B1(_0858_),
  .B2(_1533_),
  .ZN(_0345_)
);

NAND2_X1 _6371_ (
  .A1(\d_pipe[10][14] ),
  .A2(_1949_),
  .ZN(_2043_)
);

OAI21_X1 _6372_ (
  .A(_2043_),
  .B1(_0857_),
  .B2(_1944_),
  .ZN(_0346_)
);

NAND2_X1 _6373_ (
  .A1(\d_pipe[10][15] ),
  .A2(_1949_),
  .ZN(_2044_)
);

OAI21_X1 _6374_ (
  .A(_2044_),
  .B1(_0861_),
  .B2(_1944_),
  .ZN(_0347_)
);

NAND2_X1 _6375_ (
  .A1(_0926_),
  .A2(_1942_),
  .ZN(_2045_)
);

OAI21_X1 _6376_ (
  .A(_2045_),
  .B1(_0869_),
  .B2(_1944_),
  .ZN(_0348_)
);

NAND2_X1 _6377_ (
  .A1(_0931_),
  .A2(_1942_),
  .ZN(_2046_)
);

OAI21_X1 _6378_ (
  .A(_2046_),
  .B1(_0873_),
  .B2(_1944_),
  .ZN(_0349_)
);

NAND2_X1 _6379_ (
  .A1(\d_pipe[10][18] ),
  .A2(_1942_),
  .ZN(_2047_)
);

OAI21_X1 _6380_ (
  .A(_2047_),
  .B1(_0877_),
  .B2(_1944_),
  .ZN(_0350_)
);

NAND2_X1 _6381_ (
  .A1(\d_pipe[10][19] ),
  .A2(_1942_),
  .ZN(_2048_)
);

OAI21_X1 _6382_ (
  .A(_2048_),
  .B1(_0893_),
  .B2(_1535_),
  .ZN(_0351_)
);

NAND2_X1 _6383_ (
  .A1(\d_pipe[10][20] ),
  .A2(_1942_),
  .ZN(_2049_)
);

OAI21_X1 _6384_ (
  .A(_2049_),
  .B1(_0889_),
  .B2(_1535_),
  .ZN(_0352_)
);

NAND2_X1 _6385_ (
  .A1(\d_pipe[10][21] ),
  .A2(_1937_),
  .ZN(_2050_)
);

OAI21_X1 _6386_ (
  .A(_2050_),
  .B1(_0898_),
  .B2(_1535_),
  .ZN(_0353_)
);

NAND2_X1 _6387_ (
  .A1(\d_pipe[10][22] ),
  .A2(_1937_),
  .ZN(_2051_)
);

OAI21_X1 _6388_ (
  .A(_2051_),
  .B1(_0903_),
  .B2(_1535_),
  .ZN(_0354_)
);

NAND2_X1 _6389_ (
  .A1(\d_pipe[10][23] ),
  .A2(_1976_),
  .ZN(_2052_)
);

OAI21_X1 _6390_ (
  .A(_2052_),
  .B1(_0911_),
  .B2(_1539_),
  .ZN(_0355_)
);

BUF_X2 _6393_ (
  .A(_1340_),
  .Z(_2054_)
);

BUF_X1 _6399_ (
  .A(_1337_),
  .Z(_2057_)
);

MUX2_X1 _6416_ (
  .A(\s_pipe[2][2] ),
  .B(\s_pipe[1][1] ),
  .S(_1336_),
  .Z(_0368_)
);

MUX2_X1 _6417_ (
  .A(\s_pipe[2][3] ),
  .B(\s_pipe[1][2] ),
  .S(_1565_),
  .Z(_0369_)
);

BUF_X2 _6418_ (
  .A(_1346_),
  .Z(_2066_)
);

MUX2_X1 _6419_ (
  .A(\s_pipe[2][4] ),
  .B(\s_pipe[1][3] ),
  .S(_2066_),
  .Z(_0370_)
);

MUX2_X1 _6420_ (
  .A(\s_pipe[2][5] ),
  .B(\s_pipe[1][4] ),
  .S(_2066_),
  .Z(_0371_)
);

MUX2_X1 _6421_ (
  .A(\s_pipe[2][6] ),
  .B(\s_pipe[1][5] ),
  .S(_1897_),
  .Z(_0372_)
);

MUX2_X1 _6422_ (
  .A(\s_pipe[2][7] ),
  .B(\s_pipe[1][6] ),
  .S(_1898_),
  .Z(_0373_)
);

BUF_X2 _6423_ (
  .A(_1335_),
  .Z(_2067_)
);

MUX2_X1 _6424_ (
  .A(\s_pipe[2][8] ),
  .B(\s_pipe[1][7] ),
  .S(_2067_),
  .Z(_0374_)
);

MUX2_X1 _6425_ (
  .A(\s_pipe[2][9] ),
  .B(\s_pipe[1][8] ),
  .S(_2067_),
  .Z(_0375_)
);

MUX2_X1 _6426_ (
  .A(\s_pipe[2][10] ),
  .B(\s_pipe[1][9] ),
  .S(_2067_),
  .Z(_0376_)
);

BUF_X2 _6427_ (
  .A(_1335_),
  .Z(_2068_)
);

MUX2_X1 _6428_ (
  .A(\s_pipe[2][11] ),
  .B(\s_pipe[1][10] ),
  .S(_2068_),
  .Z(_0377_)
);

MUX2_X1 _6429_ (
  .A(\s_pipe[2][12] ),
  .B(_0123_),
  .S(_2068_),
  .Z(_0378_)
);

NAND2_X1 _6430_ (
  .A1(_1709_),
  .A2(\s_pipe[2][13] ),
  .ZN(_2069_)
);

OAI21_X1 _6431_ (
  .A(_2069_),
  .B1(_4060_),
  .B2(_1562_),
  .ZN(_0379_)
);

INV_X1 _6432_ (
  .A(_4059_),
  .ZN(_2070_)
);

NAND2_X1 _6433_ (
  .A1(_2070_),
  .A2(_4224_),
  .ZN(_2071_)
);

INV_X1 _6434_ (
  .A(_4224_),
  .ZN(_2072_)
);

NAND2_X1 _6435_ (
  .A1(_2072_),
  .A2(_4059_),
  .ZN(_2073_)
);

NAND3_X1 _6436_ (
  .A1(_2071_),
  .A2(_2073_),
  .A3(_1348_),
  .ZN(_2074_)
);

INV_X1 _6437_ (
  .A(\s_pipe[2][14] ),
  .ZN(_2075_)
);

OAI21_X1 _6438_ (
  .A(_2074_),
  .B1(_1408_),
  .B2(_2075_),
  .ZN(_0380_)
);

NOR2_X1 _6439_ (
  .A1(_1353_),
  .A2(\s_pipe[2][15] ),
  .ZN(_2076_)
);

INV_X1 _6440_ (
  .A(_4223_),
  .ZN(_2077_)
);

INV_X1 _6441_ (
  .A(_4220_),
  .ZN(_2078_)
);

OAI21_X2 _6442_ (
  .A(_2077_),
  .B1(_2072_),
  .B2(_2078_),
  .ZN(_2079_)
);

NAND2_X1 _6443_ (
  .A1(_4224_),
  .A2(_4221_),
  .ZN(_2080_)
);

NOR2_X1 _6444_ (
  .A1(_2080_),
  .A2(_4058_),
  .ZN(_2081_)
);

NOR2_X2 _6445_ (
  .A1(_2079_),
  .A2(_2081_),
  .ZN(_2082_)
);

INV_X1 _6446_ (
  .A(_4227_),
  .ZN(_2083_)
);

XNOR2_X1 _6447_ (
  .A(_2082_),
  .B(_2083_),
  .ZN(_2084_)
);

AOI21_X1 _6448_ (
  .A(_2076_),
  .B1(_2084_),
  .B2(_1363_),
  .ZN(_0381_)
);

NOR2_X1 _6449_ (
  .A1(_1364_),
  .A2(\s_pipe[2][16] ),
  .ZN(_2085_)
);

NOR2_X1 _6450_ (
  .A1(_4223_),
  .A2(_4226_),
  .ZN(_2086_)
);

INV_X1 _6451_ (
  .A(_4226_),
  .ZN(_2087_)
);

AOI22_X2 _6452_ (
  .A1(_2086_),
  .A2(_2071_),
  .B1(_2087_),
  .B2(_2083_),
  .ZN(_2088_)
);

BUF_X4 _6453_ (
  .A(_4230_),
  .Z(_2089_)
);

XNOR2_X1 _6454_ (
  .A(_2088_),
  .B(_2089_),
  .ZN(_2090_)
);

AOI21_X1 _6455_ (
  .A(_2085_),
  .B1(_2090_),
  .B2(_1363_),
  .ZN(_0382_)
);

BUF_X4 _6456_ (
  .A(_1347_),
  .Z(_2091_)
);

NOR2_X1 _6457_ (
  .A1(_2091_),
  .A2(\s_pipe[2][17] ),
  .ZN(_2092_)
);

INV_X1 _6458_ (
  .A(_4229_),
  .ZN(_2093_)
);

INV_X1 _6459_ (
  .A(_2089_),
  .ZN(_2094_)
);

OAI21_X1 _6460_ (
  .A(_2093_),
  .B1(_2094_),
  .B2(_2087_),
  .ZN(_2095_)
);

INV_X1 _6461_ (
  .A(_2095_),
  .ZN(_2096_)
);

NAND2_X2 _6462_ (
  .A1(_4227_),
  .A2(_2089_),
  .ZN(_2097_)
);

OAI21_X1 _6463_ (
  .A(_2096_),
  .B1(_2082_),
  .B2(_2097_),
  .ZN(_2098_)
);

BUF_X4 _6464_ (
  .A(_4233_),
  .Z(_2099_)
);

XNOR2_X1 _6465_ (
  .A(_2098_),
  .B(_2099_),
  .ZN(_2100_)
);

AOI21_X1 _6466_ (
  .A(_2092_),
  .B1(_2100_),
  .B2(_1363_),
  .ZN(_0383_)
);

NOR2_X1 _6467_ (
  .A1(_2041_),
  .A2(\s_pipe[2][18] ),
  .ZN(_2101_)
);

INV_X1 _6468_ (
  .A(_4232_),
  .ZN(_2102_)
);

INV_X1 _6469_ (
  .A(_2099_),
  .ZN(_2103_)
);

OAI21_X2 _6470_ (
  .A(_2102_),
  .B1(_2103_),
  .B2(_2093_),
  .ZN(_2104_)
);

NAND2_X1 _6471_ (
  .A1(_2089_),
  .A2(_2099_),
  .ZN(_2105_)
);

INV_X1 _6472_ (
  .A(_2105_),
  .ZN(_2106_)
);

AOI21_X1 _6473_ (
  .A(_2104_),
  .B1(_2088_),
  .B2(_2106_),
  .ZN(_2107_)
);

INV_X1 _6474_ (
  .A(_4236_),
  .ZN(_2108_)
);

XNOR2_X1 _6475_ (
  .A(_2107_),
  .B(_2108_),
  .ZN(_2109_)
);

AOI21_X1 _6476_ (
  .A(_2101_),
  .B1(_2109_),
  .B2(_1363_),
  .ZN(_0384_)
);

INV_X1 _6477_ (
  .A(_2097_),
  .ZN(_2110_)
);

NAND2_X1 _6478_ (
  .A1(_2099_),
  .A2(_4236_),
  .ZN(_2111_)
);

INV_X1 _6479_ (
  .A(_2111_),
  .ZN(_2112_)
);

NAND2_X1 _6480_ (
  .A1(_2110_),
  .A2(_2112_),
  .ZN(_2113_)
);

OR2_X2 _6481_ (
  .A1(_2082_),
  .A2(_2113_),
  .ZN(_2114_)
);

NAND2_X1 _6482_ (
  .A1(_2095_),
  .A2(_2112_),
  .ZN(_2115_)
);

INV_X1 _6483_ (
  .A(_4235_),
  .ZN(_2116_)
);

OAI21_X1 _6484_ (
  .A(_2116_),
  .B1(_2108_),
  .B2(_2102_),
  .ZN(_2117_)
);

INV_X1 _6485_ (
  .A(_2117_),
  .ZN(_2118_)
);

NAND2_X1 _6486_ (
  .A1(_2115_),
  .A2(_2118_),
  .ZN(_2119_)
);

INV_X1 _6487_ (
  .A(_2119_),
  .ZN(_2120_)
);

NAND2_X1 _6488_ (
  .A1(_2114_),
  .A2(_2120_),
  .ZN(_2121_)
);

NAND2_X1 _6489_ (
  .A1(_2121_),
  .A2(_4239_),
  .ZN(_2122_)
);

INV_X1 _6490_ (
  .A(_4239_),
  .ZN(_2123_)
);

NAND3_X1 _6491_ (
  .A1(_2114_),
  .A2(_2120_),
  .A3(_2123_),
  .ZN(_2124_)
);

NAND3_X1 _6492_ (
  .A1(_2122_),
  .A2(_2124_),
  .A3(_1348_),
  .ZN(_2125_)
);

INV_X1 _6493_ (
  .A(\s_pipe[2][19] ),
  .ZN(_2126_)
);

OAI21_X1 _6494_ (
  .A(_2125_),
  .B1(_1634_),
  .B2(_2126_),
  .ZN(_0385_)
);

NAND2_X1 _6495_ (
  .A1(_4236_),
  .A2(_4239_),
  .ZN(_2127_)
);

NOR2_X2 _6496_ (
  .A1(_2105_),
  .A2(_2127_),
  .ZN(_2128_)
);

NAND2_X1 _6497_ (
  .A1(_2088_),
  .A2(_2128_),
  .ZN(_2129_)
);

INV_X1 _6498_ (
  .A(_2127_),
  .ZN(_2130_)
);

NAND2_X1 _6499_ (
  .A1(_2104_),
  .A2(_2130_),
  .ZN(_2131_)
);

INV_X1 _6500_ (
  .A(_4238_),
  .ZN(_2132_)
);

OAI21_X1 _6501_ (
  .A(_2132_),
  .B1(_2123_),
  .B2(_2116_),
  .ZN(_2133_)
);

INV_X1 _6502_ (
  .A(_2133_),
  .ZN(_2134_)
);

NAND2_X1 _6503_ (
  .A1(_2131_),
  .A2(_2134_),
  .ZN(_2135_)
);

INV_X1 _6504_ (
  .A(_2135_),
  .ZN(_2136_)
);

NAND2_X1 _6505_ (
  .A1(_2129_),
  .A2(_2136_),
  .ZN(_2137_)
);

NAND2_X1 _6506_ (
  .A1(_2137_),
  .A2(_4242_),
  .ZN(_2138_)
);

INV_X1 _6507_ (
  .A(_4242_),
  .ZN(_2139_)
);

NAND3_X1 _6508_ (
  .A1(_2129_),
  .A2(_2136_),
  .A3(_2139_),
  .ZN(_2140_)
);

NAND3_X1 _6509_ (
  .A1(_2138_),
  .A2(_2140_),
  .A3(_1348_),
  .ZN(_2141_)
);

INV_X1 _6510_ (
  .A(\s_pipe[2][20] ),
  .ZN(_2142_)
);

OAI21_X1 _6511_ (
  .A(_2141_),
  .B1(_1901_),
  .B2(_2142_),
  .ZN(_0386_)
);

NAND2_X1 _6512_ (
  .A1(_2079_),
  .A2(_2110_),
  .ZN(_2143_)
);

NAND2_X1 _6513_ (
  .A1(_2143_),
  .A2(_2096_),
  .ZN(_2144_)
);

NAND2_X1 _6514_ (
  .A1(_4239_),
  .A2(_4242_),
  .ZN(_2145_)
);

NOR2_X1 _6515_ (
  .A1(_2111_),
  .A2(_2145_),
  .ZN(_2146_)
);

NAND2_X1 _6516_ (
  .A1(_2144_),
  .A2(_2146_),
  .ZN(_2147_)
);

INV_X1 _6517_ (
  .A(_2145_),
  .ZN(_2148_)
);

NAND2_X1 _6518_ (
  .A1(_2117_),
  .A2(_2148_),
  .ZN(_2149_)
);

INV_X1 _6519_ (
  .A(_4241_),
  .ZN(_2150_)
);

OAI21_X1 _6520_ (
  .A(_2150_),
  .B1(_2139_),
  .B2(_2132_),
  .ZN(_2151_)
);

INV_X1 _6521_ (
  .A(_2151_),
  .ZN(_2152_)
);

NAND2_X1 _6522_ (
  .A1(_2149_),
  .A2(_2152_),
  .ZN(_2153_)
);

INV_X1 _6523_ (
  .A(_2153_),
  .ZN(_2154_)
);

NOR2_X1 _6524_ (
  .A1(_2080_),
  .A2(_2097_),
  .ZN(_2155_)
);

NAND3_X1 _6525_ (
  .A1(_2155_),
  .A2(_2146_),
  .A3(_4062_),
  .ZN(_2156_)
);

NAND3_X1 _6526_ (
  .A1(_2147_),
  .A2(_2154_),
  .A3(_2156_),
  .ZN(_2157_)
);

NAND2_X1 _6527_ (
  .A1(_2157_),
  .A2(_4245_),
  .ZN(_2158_)
);

INV_X1 _6528_ (
  .A(_4245_),
  .ZN(_2159_)
);

NAND4_X1 _6529_ (
  .A1(_2147_),
  .A2(_2156_),
  .A3(_2154_),
  .A4(_2159_),
  .ZN(_2160_)
);

BUF_X2 _6530_ (
  .A(_1446_),
  .Z(_2161_)
);

NAND3_X1 _6531_ (
  .A1(_2158_),
  .A2(_2160_),
  .A3(_2161_),
  .ZN(_2162_)
);

NAND2_X1 _6532_ (
  .A1(_1490_),
  .A2(\s_pipe[2][21] ),
  .ZN(_2163_)
);

NAND2_X1 _6533_ (
  .A1(_2162_),
  .A2(_2163_),
  .ZN(_0387_)
);

OAI21_X1 _6534_ (
  .A(_2087_),
  .B1(_2083_),
  .B2(_2077_),
  .ZN(_2164_)
);

NAND2_X1 _6535_ (
  .A1(_2164_),
  .A2(_2106_),
  .ZN(_2165_)
);

INV_X1 _6536_ (
  .A(_2104_),
  .ZN(_2166_)
);

NAND2_X1 _6537_ (
  .A1(_2165_),
  .A2(_2166_),
  .ZN(_2167_)
);

NAND2_X2 _6538_ (
  .A1(_4242_),
  .A2(_4245_),
  .ZN(_2168_)
);

NOR2_X1 _6539_ (
  .A1(_2127_),
  .A2(_2168_),
  .ZN(_2169_)
);

NAND2_X1 _6540_ (
  .A1(_2167_),
  .A2(_2169_),
  .ZN(_2170_)
);

INV_X2 _6541_ (
  .A(_2168_),
  .ZN(_2171_)
);

NAND2_X1 _6542_ (
  .A1(_2133_),
  .A2(_2171_),
  .ZN(_2172_)
);

INV_X1 _6543_ (
  .A(_4244_),
  .ZN(_2173_)
);

OAI21_X1 _6544_ (
  .A(_2173_),
  .B1(_2159_),
  .B2(_2150_),
  .ZN(_2174_)
);

INV_X1 _6545_ (
  .A(_2174_),
  .ZN(_2175_)
);

NAND2_X1 _6546_ (
  .A1(_2172_),
  .A2(_2175_),
  .ZN(_2176_)
);

INV_X1 _6547_ (
  .A(_2176_),
  .ZN(_2177_)
);

NOR3_X1 _6548_ (
  .A1(_2105_),
  .A2(_2072_),
  .A3(_2083_),
  .ZN(_2178_)
);

NAND3_X1 _6549_ (
  .A1(_2178_),
  .A2(_2169_),
  .A3(_2070_),
  .ZN(_2179_)
);

NAND3_X1 _6550_ (
  .A1(_2170_),
  .A2(_2177_),
  .A3(_2179_),
  .ZN(_2180_)
);

NAND2_X1 _6551_ (
  .A1(_2180_),
  .A2(_4248_),
  .ZN(_2181_)
);

INV_X1 _6552_ (
  .A(_4248_),
  .ZN(_2182_)
);

NAND4_X1 _6553_ (
  .A1(_2170_),
  .A2(_2179_),
  .A3(_2177_),
  .A4(_2182_),
  .ZN(_2183_)
);

NAND3_X1 _6554_ (
  .A1(_2181_),
  .A2(_2183_),
  .A3(_2161_),
  .ZN(_2184_)
);

NAND2_X1 _6555_ (
  .A1(_1490_),
  .A2(\s_pipe[2][22] ),
  .ZN(_2185_)
);

NAND2_X1 _6556_ (
  .A1(_2184_),
  .A2(_2185_),
  .ZN(_0388_)
);

NAND2_X1 _6557_ (
  .A1(_4245_),
  .A2(_4248_),
  .ZN(_2186_)
);

OR2_X2 _6558_ (
  .A1(_2186_),
  .A2(_2145_),
  .ZN(_2187_)
);

INV_X1 _6559_ (
  .A(_2187_),
  .ZN(_2188_)
);

NAND2_X1 _6560_ (
  .A1(_2119_),
  .A2(_2188_),
  .ZN(_2189_)
);

INV_X1 _6561_ (
  .A(_4247_),
  .ZN(_2190_)
);

OAI21_X1 _6562_ (
  .A(_2190_),
  .B1(_2182_),
  .B2(_2173_),
  .ZN(_2191_)
);

INV_X1 _6563_ (
  .A(_2191_),
  .ZN(_2192_)
);

OAI21_X1 _6564_ (
  .A(_2192_),
  .B1(_2152_),
  .B2(_2186_),
  .ZN(_2193_)
);

INV_X1 _6565_ (
  .A(_2193_),
  .ZN(_2194_)
);

INV_X1 _6566_ (
  .A(_2082_),
  .ZN(_2195_)
);

NOR2_X2 _6567_ (
  .A1(_2187_),
  .A2(_2113_),
  .ZN(_2196_)
);

NAND2_X1 _6568_ (
  .A1(_2195_),
  .A2(_2196_),
  .ZN(_2197_)
);

INV_X1 _6569_ (
  .A(_4251_),
  .ZN(_2198_)
);

NAND4_X1 _6570_ (
  .A1(_2189_),
  .A2(_2194_),
  .A3(_2197_),
  .A4(_2198_),
  .ZN(_2199_)
);

NAND3_X1 _6571_ (
  .A1(_2189_),
  .A2(_2194_),
  .A3(_2197_),
  .ZN(_2200_)
);

NAND2_X1 _6572_ (
  .A1(_2200_),
  .A2(_4251_),
  .ZN(_2201_)
);

NAND3_X1 _6573_ (
  .A1(_2199_),
  .A2(_2201_),
  .A3(_2161_),
  .ZN(_2202_)
);

NAND2_X1 _6574_ (
  .A1(_1490_),
  .A2(\s_pipe[2][23] ),
  .ZN(_2203_)
);

NAND2_X1 _6575_ (
  .A1(_2202_),
  .A2(_2203_),
  .ZN(_0389_)
);

NAND2_X1 _6576_ (
  .A1(_4248_),
  .A2(_4251_),
  .ZN(_2204_)
);

INV_X1 _6577_ (
  .A(_2204_),
  .ZN(_2205_)
);

NAND2_X1 _6578_ (
  .A1(_2171_),
  .A2(_2205_),
  .ZN(_2206_)
);

INV_X2 _6579_ (
  .A(_2206_),
  .ZN(_2207_)
);

NAND2_X1 _6580_ (
  .A1(_2135_),
  .A2(_2207_),
  .ZN(_2208_)
);

AND2_X2 _6581_ (
  .A1(_2207_),
  .A2(_2128_),
  .ZN(_2209_)
);

NAND2_X1 _6582_ (
  .A1(_2088_),
  .A2(_2209_),
  .ZN(_2210_)
);

NAND2_X1 _6583_ (
  .A1(_2174_),
  .A2(_2205_),
  .ZN(_2211_)
);

INV_X1 _6584_ (
  .A(_4250_),
  .ZN(_2212_)
);

OAI21_X1 _6585_ (
  .A(_2212_),
  .B1(_2198_),
  .B2(_2190_),
  .ZN(_2213_)
);

INV_X1 _6586_ (
  .A(_2213_),
  .ZN(_2214_)
);

NAND2_X1 _6587_ (
  .A1(_2211_),
  .A2(_2214_),
  .ZN(_2215_)
);

INV_X1 _6588_ (
  .A(_2215_),
  .ZN(_2216_)
);

NAND3_X2 _6589_ (
  .A1(_2208_),
  .A2(_2210_),
  .A3(_2216_),
  .ZN(_2217_)
);

INV_X1 _6590_ (
  .A(_2217_),
  .ZN(_2218_)
);

NOR2_X2 _6591_ (
  .A1(_0844_),
  .A2(\d_pipe[1][23] ),
  .ZN(_2219_)
);

NAND2_X4 _6592_ (
  .A1(_0829_),
  .A2(_2219_),
  .ZN(_2220_)
);

NAND2_X2 _6593_ (
  .A1(_2220_),
  .A2(_0632_),
  .ZN(_2221_)
);

INV_X1 _6594_ (
  .A(\s_pipe[1][23] ),
  .ZN(_2222_)
);

NAND2_X1 _6595_ (
  .A1(_2221_),
  .A2(_2222_),
  .ZN(_2223_)
);

NAND3_X1 _6596_ (
  .A1(_2220_),
  .A2(_0632_),
  .A3(\s_pipe[1][23] ),
  .ZN(_2224_)
);

NAND2_X1 _6597_ (
  .A1(_2223_),
  .A2(_2224_),
  .ZN(_2225_)
);

NAND2_X1 _6598_ (
  .A1(_2218_),
  .A2(_2225_),
  .ZN(_2226_)
);

NAND2_X1 _6599_ (
  .A1(_2221_),
  .A2(\s_pipe[1][23] ),
  .ZN(_2227_)
);

NAND3_X1 _6600_ (
  .A1(_2220_),
  .A2(_0632_),
  .A3(_2222_),
  .ZN(_2228_)
);

NAND2_X1 _6601_ (
  .A1(_2227_),
  .A2(_2228_),
  .ZN(_2229_)
);

NAND2_X1 _6602_ (
  .A1(_2229_),
  .A2(_2217_),
  .ZN(_2230_)
);

NAND3_X1 _6603_ (
  .A1(_2226_),
  .A2(_2230_),
  .A3(_2161_),
  .ZN(_2231_)
);

NAND2_X1 _6604_ (
  .A1(_1449_),
  .A2(\s_pipe[2][24] ),
  .ZN(_2232_)
);

NAND2_X1 _6605_ (
  .A1(_2231_),
  .A2(_2232_),
  .ZN(_0390_)
);

MUX2_X1 _6606_ (
  .A(\s_pipe[3][3] ),
  .B(\s_pipe[2][2] ),
  .S(_1566_),
  .Z(_0391_)
);

MUX2_X1 _6607_ (
  .A(\s_pipe[3][4] ),
  .B(\s_pipe[2][3] ),
  .S(_1566_),
  .Z(_0392_)
);

MUX2_X1 _6608_ (
  .A(\s_pipe[3][5] ),
  .B(\s_pipe[2][4] ),
  .S(_1861_),
  .Z(_0393_)
);

MUX2_X1 _6609_ (
  .A(\s_pipe[3][6] ),
  .B(\s_pipe[2][5] ),
  .S(_1861_),
  .Z(_0394_)
);

MUX2_X1 _6610_ (
  .A(\s_pipe[3][7] ),
  .B(\s_pipe[2][6] ),
  .S(_1336_),
  .Z(_0395_)
);

MUX2_X1 _6611_ (
  .A(\s_pipe[3][8] ),
  .B(\s_pipe[2][7] ),
  .S(_1336_),
  .Z(_0396_)
);

MUX2_X1 _6612_ (
  .A(\s_pipe[3][9] ),
  .B(\s_pipe[2][8] ),
  .S(_1336_),
  .Z(_0397_)
);

MUX2_X1 _6613_ (
  .A(\s_pipe[3][10] ),
  .B(\s_pipe[2][9] ),
  .S(_1897_),
  .Z(_0398_)
);

MUX2_X1 _6614_ (
  .A(\s_pipe[3][11] ),
  .B(\s_pipe[2][10] ),
  .S(_1952_),
  .Z(_0399_)
);

MUX2_X1 _6615_ (
  .A(\s_pipe[3][12] ),
  .B(_0124_),
  .S(_1336_),
  .Z(_0400_)
);

NAND2_X1 _6616_ (
  .A1(_1709_),
  .A2(\s_pipe[3][13] ),
  .ZN(_2233_)
);

OAI21_X1 _6617_ (
  .A(_2233_),
  .B1(_4046_),
  .B2(_1562_),
  .ZN(_0401_)
);

INV_X1 _6618_ (
  .A(_4045_),
  .ZN(_2234_)
);

NAND2_X1 _6619_ (
  .A1(_2234_),
  .A2(_4152_),
  .ZN(_2235_)
);

INV_X1 _6620_ (
  .A(_4152_),
  .ZN(_2236_)
);

NAND2_X1 _6621_ (
  .A1(_2236_),
  .A2(_4045_),
  .ZN(_2237_)
);

BUF_X2 _6622_ (
  .A(_1347_),
  .Z(_2238_)
);

NAND3_X1 _6623_ (
  .A1(_2235_),
  .A2(_2237_),
  .A3(_2238_),
  .ZN(_2239_)
);

INV_X1 _6624_ (
  .A(\s_pipe[3][14] ),
  .ZN(_2240_)
);

OAI21_X1 _6625_ (
  .A(_2239_),
  .B1(_1408_),
  .B2(_2240_),
  .ZN(_0402_)
);

NOR2_X1 _6626_ (
  .A1(_2091_),
  .A2(\s_pipe[3][15] ),
  .ZN(_2241_)
);

INV_X1 _6627_ (
  .A(_4151_),
  .ZN(_2242_)
);

INV_X1 _6628_ (
  .A(_4148_),
  .ZN(_2243_)
);

OAI21_X2 _6629_ (
  .A(_2242_),
  .B1(_2236_),
  .B2(_2243_),
  .ZN(_2244_)
);

NAND2_X1 _6630_ (
  .A1(_4152_),
  .A2(_4149_),
  .ZN(_2245_)
);

NOR2_X1 _6631_ (
  .A1(_2245_),
  .A2(_4043_),
  .ZN(_2246_)
);

NOR2_X2 _6632_ (
  .A1(_2244_),
  .A2(_2246_),
  .ZN(_2247_)
);

INV_X1 _6633_ (
  .A(_4155_),
  .ZN(_2248_)
);

XNOR2_X1 _6634_ (
  .A(_2247_),
  .B(_2248_),
  .ZN(_2249_)
);

AOI21_X1 _6635_ (
  .A(_2241_),
  .B1(_2249_),
  .B2(_1901_),
  .ZN(_0403_)
);

NOR2_X1 _6636_ (
  .A1(_1353_),
  .A2(\s_pipe[3][16] ),
  .ZN(_2250_)
);

NOR2_X1 _6637_ (
  .A1(_4151_),
  .A2(_4154_),
  .ZN(_2251_)
);

INV_X1 _6638_ (
  .A(_4154_),
  .ZN(_2252_)
);

AOI22_X2 _6639_ (
  .A1(_2251_),
  .A2(_2235_),
  .B1(_2252_),
  .B2(_2248_),
  .ZN(_2253_)
);

BUF_X4 _6640_ (
  .A(_4158_),
  .Z(_2254_)
);

XNOR2_X1 _6641_ (
  .A(_2253_),
  .B(_2254_),
  .ZN(_2255_)
);

AOI21_X1 _6642_ (
  .A(_2250_),
  .B1(_2255_),
  .B2(_1901_),
  .ZN(_0404_)
);

NOR2_X1 _6643_ (
  .A1(_2091_),
  .A2(\s_pipe[3][17] ),
  .ZN(_2256_)
);

INV_X1 _6644_ (
  .A(_4157_),
  .ZN(_2257_)
);

INV_X1 _6645_ (
  .A(_2254_),
  .ZN(_2258_)
);

OAI21_X1 _6646_ (
  .A(_2257_),
  .B1(_2258_),
  .B2(_2252_),
  .ZN(_2259_)
);

INV_X1 _6647_ (
  .A(_2259_),
  .ZN(_2260_)
);

NAND2_X2 _6648_ (
  .A1(_4155_),
  .A2(_2254_),
  .ZN(_2261_)
);

OAI21_X1 _6649_ (
  .A(_2260_),
  .B1(_2247_),
  .B2(_2261_),
  .ZN(_2262_)
);

BUF_X4 _6650_ (
  .A(_4161_),
  .Z(_2263_)
);

XNOR2_X1 _6651_ (
  .A(_2262_),
  .B(_2263_),
  .ZN(_2264_)
);

BUF_X2 _6652_ (
  .A(_1350_),
  .Z(_2265_)
);

AOI21_X1 _6653_ (
  .A(_2256_),
  .B1(_2264_),
  .B2(_2265_),
  .ZN(_0405_)
);

NOR2_X1 _6654_ (
  .A1(_1371_),
  .A2(\s_pipe[3][18] ),
  .ZN(_2266_)
);

INV_X1 _6655_ (
  .A(_4160_),
  .ZN(_2267_)
);

INV_X1 _6656_ (
  .A(_2263_),
  .ZN(_2268_)
);

OAI21_X2 _6657_ (
  .A(_2267_),
  .B1(_2268_),
  .B2(_2257_),
  .ZN(_2269_)
);

NAND2_X1 _6658_ (
  .A1(_2254_),
  .A2(_2263_),
  .ZN(_2270_)
);

INV_X1 _6659_ (
  .A(_2270_),
  .ZN(_2271_)
);

AOI21_X1 _6660_ (
  .A(_2269_),
  .B1(_2253_),
  .B2(_2271_),
  .ZN(_2272_)
);

INV_X1 _6661_ (
  .A(_4164_),
  .ZN(_2273_)
);

XNOR2_X1 _6662_ (
  .A(_2272_),
  .B(_2273_),
  .ZN(_2274_)
);

AOI21_X1 _6663_ (
  .A(_2266_),
  .B1(_2274_),
  .B2(_2265_),
  .ZN(_0406_)
);

INV_X1 _6664_ (
  .A(_2261_),
  .ZN(_2275_)
);

NAND2_X1 _6665_ (
  .A1(_2263_),
  .A2(_4164_),
  .ZN(_2276_)
);

INV_X1 _6666_ (
  .A(_2276_),
  .ZN(_2277_)
);

NAND2_X1 _6667_ (
  .A1(_2275_),
  .A2(_2277_),
  .ZN(_2278_)
);

OR2_X2 _6668_ (
  .A1(_2247_),
  .A2(_2278_),
  .ZN(_2279_)
);

NAND2_X1 _6669_ (
  .A1(_2259_),
  .A2(_2277_),
  .ZN(_2280_)
);

INV_X1 _6670_ (
  .A(_4163_),
  .ZN(_2281_)
);

OAI21_X1 _6671_ (
  .A(_2281_),
  .B1(_2273_),
  .B2(_2267_),
  .ZN(_2282_)
);

INV_X1 _6672_ (
  .A(_2282_),
  .ZN(_2283_)
);

NAND2_X1 _6673_ (
  .A1(_2280_),
  .A2(_2283_),
  .ZN(_2284_)
);

INV_X1 _6674_ (
  .A(_2284_),
  .ZN(_2285_)
);

NAND2_X1 _6675_ (
  .A1(_2279_),
  .A2(_2285_),
  .ZN(_2286_)
);

NAND2_X1 _6676_ (
  .A1(_2286_),
  .A2(_4167_),
  .ZN(_2287_)
);

INV_X1 _6677_ (
  .A(_4167_),
  .ZN(_2288_)
);

NAND3_X1 _6678_ (
  .A1(_2279_),
  .A2(_2285_),
  .A3(_2288_),
  .ZN(_2289_)
);

NAND3_X1 _6679_ (
  .A1(_2287_),
  .A2(_2289_),
  .A3(_2238_),
  .ZN(_2290_)
);

BUF_X2 _6680_ (
  .A(_1350_),
  .Z(_2291_)
);

INV_X1 _6681_ (
  .A(\s_pipe[3][19] ),
  .ZN(_2292_)
);

OAI21_X1 _6682_ (
  .A(_2290_),
  .B1(_2291_),
  .B2(_2292_),
  .ZN(_0407_)
);

NAND2_X1 _6683_ (
  .A1(_4164_),
  .A2(_4167_),
  .ZN(_2293_)
);

NOR2_X2 _6684_ (
  .A1(_2270_),
  .A2(_2293_),
  .ZN(_2294_)
);

NAND2_X1 _6685_ (
  .A1(_2253_),
  .A2(_2294_),
  .ZN(_2295_)
);

INV_X1 _6686_ (
  .A(_2293_),
  .ZN(_2296_)
);

NAND2_X1 _6687_ (
  .A1(_2269_),
  .A2(_2296_),
  .ZN(_2297_)
);

INV_X1 _6688_ (
  .A(_4166_),
  .ZN(_2298_)
);

OAI21_X1 _6689_ (
  .A(_2298_),
  .B1(_2288_),
  .B2(_2281_),
  .ZN(_2299_)
);

INV_X1 _6690_ (
  .A(_2299_),
  .ZN(_2300_)
);

NAND2_X1 _6691_ (
  .A1(_2297_),
  .A2(_2300_),
  .ZN(_2301_)
);

INV_X1 _6692_ (
  .A(_2301_),
  .ZN(_2302_)
);

NAND2_X1 _6693_ (
  .A1(_2295_),
  .A2(_2302_),
  .ZN(_2303_)
);

NAND2_X1 _6694_ (
  .A1(_2303_),
  .A2(_4170_),
  .ZN(_2304_)
);

INV_X1 _6695_ (
  .A(_4170_),
  .ZN(_2305_)
);

NAND3_X1 _6696_ (
  .A1(_2295_),
  .A2(_2302_),
  .A3(_2305_),
  .ZN(_2306_)
);

NAND3_X1 _6697_ (
  .A1(_2304_),
  .A2(_2306_),
  .A3(_2238_),
  .ZN(_2307_)
);

INV_X1 _6698_ (
  .A(\s_pipe[3][20] ),
  .ZN(_2308_)
);

OAI21_X1 _6699_ (
  .A(_2307_),
  .B1(_2291_),
  .B2(_2308_),
  .ZN(_0408_)
);

NAND2_X1 _6700_ (
  .A1(_2244_),
  .A2(_2275_),
  .ZN(_2309_)
);

NAND2_X1 _6701_ (
  .A1(_2309_),
  .A2(_2260_),
  .ZN(_2310_)
);

NAND2_X1 _6702_ (
  .A1(_4167_),
  .A2(_4170_),
  .ZN(_2311_)
);

NOR2_X1 _6703_ (
  .A1(_2276_),
  .A2(_2311_),
  .ZN(_2312_)
);

NAND2_X1 _6704_ (
  .A1(_2310_),
  .A2(_2312_),
  .ZN(_2313_)
);

INV_X1 _6705_ (
  .A(_2311_),
  .ZN(_2314_)
);

NAND2_X1 _6706_ (
  .A1(_2282_),
  .A2(_2314_),
  .ZN(_2315_)
);

INV_X1 _6707_ (
  .A(_4169_),
  .ZN(_2316_)
);

OAI21_X1 _6708_ (
  .A(_2316_),
  .B1(_2305_),
  .B2(_2298_),
  .ZN(_2317_)
);

INV_X1 _6709_ (
  .A(_2317_),
  .ZN(_2318_)
);

NAND2_X1 _6710_ (
  .A1(_2315_),
  .A2(_2318_),
  .ZN(_2319_)
);

INV_X1 _6711_ (
  .A(_2319_),
  .ZN(_2320_)
);

NOR2_X1 _6712_ (
  .A1(_2245_),
  .A2(_2261_),
  .ZN(_2321_)
);

NAND3_X1 _6713_ (
  .A1(_2321_),
  .A2(_2312_),
  .A3(_4047_),
  .ZN(_2322_)
);

NAND3_X1 _6714_ (
  .A1(_2313_),
  .A2(_2320_),
  .A3(_2322_),
  .ZN(_2323_)
);

NAND2_X1 _6715_ (
  .A1(_2323_),
  .A2(_4173_),
  .ZN(_2324_)
);

INV_X1 _6716_ (
  .A(_4173_),
  .ZN(_2325_)
);

NAND4_X1 _6717_ (
  .A1(_2313_),
  .A2(_2322_),
  .A3(_2320_),
  .A4(_2325_),
  .ZN(_2326_)
);

NAND3_X1 _6718_ (
  .A1(_2324_),
  .A2(_2326_),
  .A3(_2001_),
  .ZN(_2327_)
);

NAND2_X1 _6719_ (
  .A1(_1449_),
  .A2(\s_pipe[3][21] ),
  .ZN(_2328_)
);

NAND2_X1 _6720_ (
  .A1(_2327_),
  .A2(_2328_),
  .ZN(_0409_)
);

OAI21_X1 _6721_ (
  .A(_2252_),
  .B1(_2248_),
  .B2(_2242_),
  .ZN(_2329_)
);

NAND2_X1 _6722_ (
  .A1(_2329_),
  .A2(_2271_),
  .ZN(_2330_)
);

INV_X1 _6723_ (
  .A(_2269_),
  .ZN(_2331_)
);

NAND2_X1 _6724_ (
  .A1(_2330_),
  .A2(_2331_),
  .ZN(_2332_)
);

NAND2_X1 _6725_ (
  .A1(_4170_),
  .A2(_4173_),
  .ZN(_2333_)
);

NOR2_X1 _6726_ (
  .A1(_2293_),
  .A2(_2333_),
  .ZN(_2334_)
);

NAND2_X1 _6727_ (
  .A1(_2332_),
  .A2(_2334_),
  .ZN(_2335_)
);

INV_X2 _6728_ (
  .A(_2333_),
  .ZN(_2336_)
);

NAND2_X1 _6729_ (
  .A1(_2299_),
  .A2(_2336_),
  .ZN(_2337_)
);

INV_X1 _6730_ (
  .A(_4172_),
  .ZN(_2338_)
);

OAI21_X1 _6731_ (
  .A(_2338_),
  .B1(_2325_),
  .B2(_2316_),
  .ZN(_2339_)
);

INV_X1 _6732_ (
  .A(_2339_),
  .ZN(_2340_)
);

NAND2_X1 _6733_ (
  .A1(_2337_),
  .A2(_2340_),
  .ZN(_2341_)
);

INV_X1 _6734_ (
  .A(_2341_),
  .ZN(_2342_)
);

NOR3_X1 _6735_ (
  .A1(_2270_),
  .A2(_2236_),
  .A3(_2248_),
  .ZN(_2343_)
);

NAND3_X1 _6736_ (
  .A1(_2343_),
  .A2(_2334_),
  .A3(_2234_),
  .ZN(_2344_)
);

NAND3_X1 _6737_ (
  .A1(_2335_),
  .A2(_2342_),
  .A3(_2344_),
  .ZN(_2345_)
);

NAND2_X1 _6738_ (
  .A1(_2345_),
  .A2(_4176_),
  .ZN(_2346_)
);

INV_X1 _6739_ (
  .A(_4176_),
  .ZN(_2347_)
);

NAND4_X1 _6740_ (
  .A1(_2335_),
  .A2(_2344_),
  .A3(_2342_),
  .A4(_2347_),
  .ZN(_2348_)
);

BUF_X2 _6741_ (
  .A(_1446_),
  .Z(_2349_)
);

NAND3_X1 _6742_ (
  .A1(_2346_),
  .A2(_2348_),
  .A3(_2349_),
  .ZN(_2350_)
);

NAND2_X1 _6743_ (
  .A1(_1449_),
  .A2(\s_pipe[3][22] ),
  .ZN(_2351_)
);

NAND2_X1 _6744_ (
  .A1(_2350_),
  .A2(_2351_),
  .ZN(_0410_)
);

NAND2_X1 _6745_ (
  .A1(_4173_),
  .A2(_4176_),
  .ZN(_2352_)
);

OR2_X2 _6746_ (
  .A1(_2352_),
  .A2(_2311_),
  .ZN(_2353_)
);

INV_X1 _6747_ (
  .A(_2353_),
  .ZN(_2354_)
);

NAND2_X1 _6748_ (
  .A1(_2284_),
  .A2(_2354_),
  .ZN(_2355_)
);

INV_X1 _6749_ (
  .A(_4175_),
  .ZN(_2356_)
);

OAI21_X1 _6750_ (
  .A(_2356_),
  .B1(_2347_),
  .B2(_2338_),
  .ZN(_2357_)
);

INV_X1 _6751_ (
  .A(_2357_),
  .ZN(_2358_)
);

OAI21_X1 _6752_ (
  .A(_2358_),
  .B1(_2318_),
  .B2(_2352_),
  .ZN(_2359_)
);

INV_X1 _6753_ (
  .A(_2359_),
  .ZN(_2360_)
);

INV_X1 _6754_ (
  .A(_2247_),
  .ZN(_2361_)
);

NOR2_X2 _6755_ (
  .A1(_2353_),
  .A2(_2278_),
  .ZN(_2362_)
);

NAND2_X1 _6756_ (
  .A1(_2361_),
  .A2(_2362_),
  .ZN(_2363_)
);

INV_X1 _6757_ (
  .A(_4179_),
  .ZN(_2364_)
);

NAND4_X1 _6758_ (
  .A1(_2355_),
  .A2(_2360_),
  .A3(_2363_),
  .A4(_2364_),
  .ZN(_2365_)
);

NAND3_X1 _6759_ (
  .A1(_2355_),
  .A2(_2360_),
  .A3(_2363_),
  .ZN(_2366_)
);

NAND2_X1 _6760_ (
  .A1(_2366_),
  .A2(_4179_),
  .ZN(_2367_)
);

NAND3_X1 _6761_ (
  .A1(_2365_),
  .A2(_2367_),
  .A3(_2349_),
  .ZN(_2368_)
);

NAND2_X1 _6762_ (
  .A1(_1449_),
  .A2(\s_pipe[3][23] ),
  .ZN(_2369_)
);

NAND2_X1 _6763_ (
  .A1(_2368_),
  .A2(_2369_),
  .ZN(_0411_)
);

NAND2_X1 _6764_ (
  .A1(_4176_),
  .A2(_4179_),
  .ZN(_2370_)
);

INV_X1 _6765_ (
  .A(_2370_),
  .ZN(_2371_)
);

NAND2_X1 _6766_ (
  .A1(_2336_),
  .A2(_2371_),
  .ZN(_2372_)
);

INV_X2 _6767_ (
  .A(_2372_),
  .ZN(_2373_)
);

NAND2_X1 _6768_ (
  .A1(_2301_),
  .A2(_2373_),
  .ZN(_2374_)
);

AND2_X2 _6769_ (
  .A1(_2373_),
  .A2(_2294_),
  .ZN(_2375_)
);

NAND2_X2 _6770_ (
  .A1(_2253_),
  .A2(_2375_),
  .ZN(_2376_)
);

NAND2_X1 _6771_ (
  .A1(_2339_),
  .A2(_2371_),
  .ZN(_2377_)
);

INV_X1 _6772_ (
  .A(_4178_),
  .ZN(_2378_)
);

OAI21_X1 _6773_ (
  .A(_2378_),
  .B1(_2364_),
  .B2(_2356_),
  .ZN(_2379_)
);

INV_X1 _6774_ (
  .A(_2379_),
  .ZN(_2380_)
);

NAND2_X1 _6775_ (
  .A1(_2377_),
  .A2(_2380_),
  .ZN(_2381_)
);

INV_X1 _6776_ (
  .A(_2381_),
  .ZN(_2382_)
);

NAND3_X2 _6777_ (
  .A1(_2374_),
  .A2(_2376_),
  .A3(_2382_),
  .ZN(_2383_)
);

INV_X1 _6778_ (
  .A(_2383_),
  .ZN(_2384_)
);

NOR2_X2 _6779_ (
  .A1(_0731_),
  .A2(_0738_),
  .ZN(_2385_)
);

NAND2_X4 _6780_ (
  .A1(_0714_),
  .A2(_2385_),
  .ZN(_2386_)
);

NAND2_X4 _6781_ (
  .A1(_2386_),
  .A2(_0626_),
  .ZN(_2387_)
);

INV_X1 _6782_ (
  .A(\s_pipe[2][23] ),
  .ZN(_2388_)
);

NAND2_X1 _6783_ (
  .A1(_2387_),
  .A2(_2388_),
  .ZN(_2389_)
);

NAND3_X1 _6784_ (
  .A1(_2386_),
  .A2(_0626_),
  .A3(\s_pipe[2][23] ),
  .ZN(_2390_)
);

NAND2_X1 _6785_ (
  .A1(_2389_),
  .A2(_2390_),
  .ZN(_2391_)
);

NAND2_X1 _6786_ (
  .A1(_2384_),
  .A2(_2391_),
  .ZN(_2392_)
);

NAND2_X1 _6787_ (
  .A1(_2387_),
  .A2(\s_pipe[2][23] ),
  .ZN(_2393_)
);

NAND3_X1 _6788_ (
  .A1(_2386_),
  .A2(_0626_),
  .A3(_2388_),
  .ZN(_2394_)
);

NAND2_X1 _6789_ (
  .A1(_2393_),
  .A2(_2394_),
  .ZN(_2395_)
);

NAND2_X1 _6790_ (
  .A1(_2395_),
  .A2(_2383_),
  .ZN(_2396_)
);

NAND3_X1 _6791_ (
  .A1(_2392_),
  .A2(_2396_),
  .A3(_2349_),
  .ZN(_2397_)
);

NAND2_X1 _6792_ (
  .A1(_1449_),
  .A2(\s_pipe[3][24] ),
  .ZN(_2398_)
);

NAND2_X1 _6793_ (
  .A1(_2397_),
  .A2(_2398_),
  .ZN(_0412_)
);

NAND2_X1 _6794_ (
  .A1(_1709_),
  .A2(\s_pipe[11][11] ),
  .ZN(_2399_)
);

INV_X1 _6795_ (
  .A(\s_pipe[10][10] ),
  .ZN(_2400_)
);

OAI21_X1 _6796_ (
  .A(_2399_),
  .B1(_1524_),
  .B2(_2400_),
  .ZN(_0413_)
);

MUX2_X1 _6797_ (
  .A(\s_pipe[11][12] ),
  .B(_0141_),
  .S(_2007_),
  .Z(_0414_)
);

NAND2_X1 _6798_ (
  .A1(_1881_),
  .A2(\s_pipe[11][13] ),
  .ZN(_2401_)
);

OAI21_X1 _6799_ (
  .A(_2401_),
  .B1(_4077_),
  .B2(_1341_),
  .ZN(_0415_)
);

INV_X1 _6800_ (
  .A(_4076_),
  .ZN(_2402_)
);

NAND2_X1 _6801_ (
  .A1(_2402_),
  .A2(_4329_),
  .ZN(_2403_)
);

INV_X1 _6802_ (
  .A(_4329_),
  .ZN(_2404_)
);

NAND2_X1 _6803_ (
  .A1(_2404_),
  .A2(_4076_),
  .ZN(_2405_)
);

NAND3_X1 _6804_ (
  .A1(_2403_),
  .A2(_2405_),
  .A3(_2238_),
  .ZN(_2406_)
);

INV_X1 _6805_ (
  .A(\s_pipe[11][14] ),
  .ZN(_2407_)
);

OAI21_X1 _6806_ (
  .A(_2406_),
  .B1(_2291_),
  .B2(_2407_),
  .ZN(_0416_)
);

NOR2_X1 _6807_ (
  .A1(_2091_),
  .A2(\s_pipe[11][15] ),
  .ZN(_2408_)
);

INV_X1 _6808_ (
  .A(_4328_),
  .ZN(_2409_)
);

INV_X1 _6809_ (
  .A(_4325_),
  .ZN(_2410_)
);

OAI21_X2 _6810_ (
  .A(_2409_),
  .B1(_2404_),
  .B2(_2410_),
  .ZN(_2411_)
);

NAND2_X1 _6811_ (
  .A1(_4329_),
  .A2(_4326_),
  .ZN(_2412_)
);

NOR2_X1 _6812_ (
  .A1(_2412_),
  .A2(_4075_),
  .ZN(_2413_)
);

NOR2_X2 _6813_ (
  .A1(_2411_),
  .A2(_2413_),
  .ZN(_2414_)
);

INV_X1 _6814_ (
  .A(_4332_),
  .ZN(_2415_)
);

XNOR2_X1 _6815_ (
  .A(_2414_),
  .B(_2415_),
  .ZN(_2416_)
);

AOI21_X1 _6816_ (
  .A(_2408_),
  .B1(_2416_),
  .B2(_1587_),
  .ZN(_0417_)
);

NOR2_X1 _6817_ (
  .A1(_2091_),
  .A2(\s_pipe[11][16] ),
  .ZN(_2417_)
);

NOR2_X1 _6818_ (
  .A1(_4328_),
  .A2(_4331_),
  .ZN(_2418_)
);

INV_X1 _6819_ (
  .A(_4331_),
  .ZN(_2419_)
);

AOI22_X2 _6820_ (
  .A1(_2418_),
  .A2(_2403_),
  .B1(_2419_),
  .B2(_2415_),
  .ZN(_2420_)
);

BUF_X4 _6821_ (
  .A(_4335_),
  .Z(_2421_)
);

XNOR2_X1 _6822_ (
  .A(_2420_),
  .B(_2421_),
  .ZN(_2422_)
);

AOI21_X1 _6823_ (
  .A(_2417_),
  .B1(_2422_),
  .B2(_1587_),
  .ZN(_0418_)
);

NOR2_X1 _6824_ (
  .A1(_2091_),
  .A2(\s_pipe[11][17] ),
  .ZN(_2423_)
);

INV_X1 _6825_ (
  .A(_4334_),
  .ZN(_2424_)
);

INV_X1 _6826_ (
  .A(_2421_),
  .ZN(_2425_)
);

OAI21_X1 _6827_ (
  .A(_2424_),
  .B1(_2425_),
  .B2(_2419_),
  .ZN(_2426_)
);

INV_X1 _6828_ (
  .A(_2426_),
  .ZN(_2427_)
);

NAND2_X2 _6829_ (
  .A1(_4332_),
  .A2(_2421_),
  .ZN(_2428_)
);

OAI21_X1 _6830_ (
  .A(_2427_),
  .B1(_2414_),
  .B2(_2428_),
  .ZN(_2429_)
);

BUF_X4 _6831_ (
  .A(_4338_),
  .Z(_2430_)
);

XNOR2_X1 _6832_ (
  .A(_2429_),
  .B(_2430_),
  .ZN(_2431_)
);

AOI21_X1 _6833_ (
  .A(_2423_),
  .B1(_2431_),
  .B2(_1363_),
  .ZN(_0419_)
);

NOR2_X1 _6834_ (
  .A1(_1364_),
  .A2(\s_pipe[11][18] ),
  .ZN(_2432_)
);

INV_X1 _6835_ (
  .A(_4337_),
  .ZN(_2433_)
);

INV_X1 _6836_ (
  .A(_2430_),
  .ZN(_2434_)
);

OAI21_X2 _6837_ (
  .A(_2433_),
  .B1(_2434_),
  .B2(_2424_),
  .ZN(_2435_)
);

NAND2_X1 _6838_ (
  .A1(_2421_),
  .A2(_2430_),
  .ZN(_2436_)
);

INV_X1 _6839_ (
  .A(_2436_),
  .ZN(_2437_)
);

AOI21_X1 _6840_ (
  .A(_2435_),
  .B1(_2420_),
  .B2(_2437_),
  .ZN(_2438_)
);

INV_X1 _6841_ (
  .A(_4341_),
  .ZN(_2439_)
);

XNOR2_X1 _6842_ (
  .A(_2438_),
  .B(_2439_),
  .ZN(_2440_)
);

AOI21_X1 _6843_ (
  .A(_2432_),
  .B1(_2440_),
  .B2(_1381_),
  .ZN(_0420_)
);

INV_X1 _6844_ (
  .A(_2428_),
  .ZN(_2441_)
);

NAND2_X1 _6845_ (
  .A1(_2430_),
  .A2(_4341_),
  .ZN(_2442_)
);

INV_X1 _6846_ (
  .A(_2442_),
  .ZN(_2443_)
);

NAND2_X1 _6847_ (
  .A1(_2441_),
  .A2(_2443_),
  .ZN(_2444_)
);

OR2_X2 _6848_ (
  .A1(_2414_),
  .A2(_2444_),
  .ZN(_2445_)
);

NAND2_X1 _6849_ (
  .A1(_2426_),
  .A2(_2443_),
  .ZN(_2446_)
);

INV_X1 _6850_ (
  .A(_4340_),
  .ZN(_2447_)
);

OAI21_X1 _6851_ (
  .A(_2447_),
  .B1(_2439_),
  .B2(_2433_),
  .ZN(_2448_)
);

INV_X1 _6852_ (
  .A(_2448_),
  .ZN(_2449_)
);

NAND2_X1 _6853_ (
  .A1(_2446_),
  .A2(_2449_),
  .ZN(_2450_)
);

INV_X1 _6854_ (
  .A(_2450_),
  .ZN(_2451_)
);

NAND2_X1 _6855_ (
  .A1(_2445_),
  .A2(_2451_),
  .ZN(_2452_)
);

NAND2_X1 _6856_ (
  .A1(_2452_),
  .A2(_4344_),
  .ZN(_2453_)
);

INV_X1 _6857_ (
  .A(_4344_),
  .ZN(_2454_)
);

NAND3_X1 _6858_ (
  .A1(_2445_),
  .A2(_2451_),
  .A3(_2454_),
  .ZN(_2455_)
);

NAND3_X1 _6859_ (
  .A1(_2453_),
  .A2(_2455_),
  .A3(_1572_),
  .ZN(_2456_)
);

INV_X1 _6860_ (
  .A(\s_pipe[11][19] ),
  .ZN(_2457_)
);

OAI21_X1 _6861_ (
  .A(_2456_),
  .B1(_1408_),
  .B2(_2457_),
  .ZN(_0421_)
);

NAND2_X1 _6862_ (
  .A1(_4341_),
  .A2(_4344_),
  .ZN(_2458_)
);

NOR2_X2 _6863_ (
  .A1(_2436_),
  .A2(_2458_),
  .ZN(_2459_)
);

NAND2_X1 _6864_ (
  .A1(_2420_),
  .A2(_2459_),
  .ZN(_2460_)
);

INV_X1 _6865_ (
  .A(_2458_),
  .ZN(_2461_)
);

NAND2_X1 _6866_ (
  .A1(_2435_),
  .A2(_2461_),
  .ZN(_2462_)
);

INV_X1 _6867_ (
  .A(_4343_),
  .ZN(_2463_)
);

OAI21_X1 _6868_ (
  .A(_2463_),
  .B1(_2454_),
  .B2(_2447_),
  .ZN(_2464_)
);

INV_X1 _6869_ (
  .A(_2464_),
  .ZN(_2465_)
);

NAND2_X1 _6870_ (
  .A1(_2462_),
  .A2(_2465_),
  .ZN(_2466_)
);

INV_X1 _6871_ (
  .A(_2466_),
  .ZN(_2467_)
);

NAND2_X1 _6872_ (
  .A1(_2460_),
  .A2(_2467_),
  .ZN(_2468_)
);

NAND2_X1 _6873_ (
  .A1(_2468_),
  .A2(_4347_),
  .ZN(_2469_)
);

INV_X1 _6874_ (
  .A(_4347_),
  .ZN(_2470_)
);

NAND3_X1 _6875_ (
  .A1(_2460_),
  .A2(_2467_),
  .A3(_2470_),
  .ZN(_2471_)
);

NAND3_X1 _6876_ (
  .A1(_2469_),
  .A2(_2471_),
  .A3(_1572_),
  .ZN(_2472_)
);

INV_X1 _6877_ (
  .A(\s_pipe[11][20] ),
  .ZN(_2473_)
);

OAI21_X1 _6878_ (
  .A(_2472_),
  .B1(_1408_),
  .B2(_2473_),
  .ZN(_0422_)
);

NAND2_X1 _6879_ (
  .A1(_2411_),
  .A2(_2441_),
  .ZN(_2474_)
);

NAND2_X1 _6880_ (
  .A1(_2474_),
  .A2(_2427_),
  .ZN(_2475_)
);

NAND2_X1 _6881_ (
  .A1(_4344_),
  .A2(_4347_),
  .ZN(_2476_)
);

NOR2_X1 _6882_ (
  .A1(_2442_),
  .A2(_2476_),
  .ZN(_2477_)
);

NAND2_X1 _6883_ (
  .A1(_2475_),
  .A2(_2477_),
  .ZN(_2478_)
);

INV_X1 _6884_ (
  .A(_2476_),
  .ZN(_2479_)
);

NAND2_X1 _6885_ (
  .A1(_2448_),
  .A2(_2479_),
  .ZN(_2480_)
);

INV_X1 _6886_ (
  .A(_4346_),
  .ZN(_2481_)
);

OAI21_X1 _6887_ (
  .A(_2481_),
  .B1(_2470_),
  .B2(_2463_),
  .ZN(_2482_)
);

INV_X1 _6888_ (
  .A(_2482_),
  .ZN(_2483_)
);

NAND2_X1 _6889_ (
  .A1(_2480_),
  .A2(_2483_),
  .ZN(_2484_)
);

INV_X1 _6890_ (
  .A(_2484_),
  .ZN(_2485_)
);

NOR2_X1 _6891_ (
  .A1(_2412_),
  .A2(_2428_),
  .ZN(_2486_)
);

NAND3_X1 _6892_ (
  .A1(_2486_),
  .A2(_2477_),
  .A3(_4079_),
  .ZN(_2487_)
);

NAND3_X1 _6893_ (
  .A1(_2478_),
  .A2(_2485_),
  .A3(_2487_),
  .ZN(_2488_)
);

NAND2_X1 _6894_ (
  .A1(_2488_),
  .A2(_4350_),
  .ZN(_2489_)
);

INV_X1 _6895_ (
  .A(_4350_),
  .ZN(_2490_)
);

NAND4_X1 _6896_ (
  .A1(_2478_),
  .A2(_2487_),
  .A3(_2485_),
  .A4(_2490_),
  .ZN(_2491_)
);

NAND3_X1 _6897_ (
  .A1(_2489_),
  .A2(_2491_),
  .A3(_1447_),
  .ZN(_2492_)
);

NAND2_X1 _6898_ (
  .A1(_1341_),
  .A2(\s_pipe[11][21] ),
  .ZN(_2493_)
);

NAND2_X1 _6899_ (
  .A1(_2492_),
  .A2(_2493_),
  .ZN(_0423_)
);

OAI21_X1 _6900_ (
  .A(_2419_),
  .B1(_2415_),
  .B2(_2409_),
  .ZN(_2494_)
);

NAND2_X1 _6901_ (
  .A1(_2494_),
  .A2(_2437_),
  .ZN(_2495_)
);

INV_X1 _6902_ (
  .A(_2435_),
  .ZN(_2496_)
);

NAND2_X1 _6903_ (
  .A1(_2495_),
  .A2(_2496_),
  .ZN(_2497_)
);

NAND2_X1 _6904_ (
  .A1(_4347_),
  .A2(_4350_),
  .ZN(_2498_)
);

NOR2_X1 _6905_ (
  .A1(_2458_),
  .A2(_2498_),
  .ZN(_2499_)
);

NAND2_X1 _6906_ (
  .A1(_2497_),
  .A2(_2499_),
  .ZN(_2500_)
);

INV_X2 _6907_ (
  .A(_2498_),
  .ZN(_2501_)
);

NAND2_X1 _6908_ (
  .A1(_2464_),
  .A2(_2501_),
  .ZN(_2502_)
);

INV_X1 _6909_ (
  .A(_4349_),
  .ZN(_2503_)
);

OAI21_X1 _6910_ (
  .A(_2503_),
  .B1(_2490_),
  .B2(_2481_),
  .ZN(_2504_)
);

INV_X1 _6911_ (
  .A(_2504_),
  .ZN(_2505_)
);

NAND2_X1 _6912_ (
  .A1(_2502_),
  .A2(_2505_),
  .ZN(_2506_)
);

INV_X1 _6913_ (
  .A(_2506_),
  .ZN(_2507_)
);

NOR3_X1 _6914_ (
  .A1(_2436_),
  .A2(_2404_),
  .A3(_2415_),
  .ZN(_2508_)
);

NAND3_X1 _6915_ (
  .A1(_2508_),
  .A2(_2499_),
  .A3(_2402_),
  .ZN(_2509_)
);

NAND3_X1 _6916_ (
  .A1(_2500_),
  .A2(_2507_),
  .A3(_2509_),
  .ZN(_2510_)
);

NAND2_X1 _6917_ (
  .A1(_2510_),
  .A2(_4353_),
  .ZN(_2511_)
);

INV_X1 _6918_ (
  .A(_4353_),
  .ZN(_2512_)
);

NAND4_X1 _6919_ (
  .A1(_2500_),
  .A2(_2509_),
  .A3(_2507_),
  .A4(_2512_),
  .ZN(_2513_)
);

NAND3_X1 _6920_ (
  .A1(_2511_),
  .A2(_2513_),
  .A3(_2001_),
  .ZN(_2514_)
);

NAND2_X1 _6921_ (
  .A1(_1449_),
  .A2(\s_pipe[11][22] ),
  .ZN(_2515_)
);

NAND2_X1 _6922_ (
  .A1(_2514_),
  .A2(_2515_),
  .ZN(_0424_)
);

NAND2_X1 _6923_ (
  .A1(_4350_),
  .A2(_4353_),
  .ZN(_2516_)
);

OR2_X2 _6924_ (
  .A1(_2516_),
  .A2(_2476_),
  .ZN(_2517_)
);

INV_X1 _6925_ (
  .A(_2517_),
  .ZN(_2518_)
);

NAND2_X1 _6926_ (
  .A1(_2450_),
  .A2(_2518_),
  .ZN(_2519_)
);

INV_X1 _6927_ (
  .A(_4352_),
  .ZN(_2520_)
);

OAI21_X1 _6928_ (
  .A(_2520_),
  .B1(_2512_),
  .B2(_2503_),
  .ZN(_2521_)
);

INV_X1 _6929_ (
  .A(_2521_),
  .ZN(_2522_)
);

OAI21_X1 _6930_ (
  .A(_2522_),
  .B1(_2483_),
  .B2(_2516_),
  .ZN(_2523_)
);

INV_X1 _6931_ (
  .A(_2523_),
  .ZN(_2524_)
);

INV_X1 _6932_ (
  .A(_2414_),
  .ZN(_2525_)
);

NOR2_X2 _6933_ (
  .A1(_2517_),
  .A2(_2444_),
  .ZN(_2526_)
);

NAND2_X1 _6934_ (
  .A1(_2525_),
  .A2(_2526_),
  .ZN(_2527_)
);

INV_X1 _6935_ (
  .A(_4356_),
  .ZN(_2528_)
);

NAND4_X1 _6936_ (
  .A1(_2519_),
  .A2(_2524_),
  .A3(_2527_),
  .A4(_2528_),
  .ZN(_2529_)
);

NAND3_X1 _6937_ (
  .A1(_2519_),
  .A2(_2524_),
  .A3(_2527_),
  .ZN(_2530_)
);

NAND2_X1 _6938_ (
  .A1(_2530_),
  .A2(_4356_),
  .ZN(_2531_)
);

NAND3_X1 _6939_ (
  .A1(_2529_),
  .A2(_2531_),
  .A3(_1447_),
  .ZN(_2532_)
);

NAND2_X1 _6940_ (
  .A1(_1709_),
  .A2(\s_pipe[11][23] ),
  .ZN(_2533_)
);

NAND2_X1 _6941_ (
  .A1(_2532_),
  .A2(_2533_),
  .ZN(_0425_)
);

NAND2_X1 _6942_ (
  .A1(_4353_),
  .A2(_4356_),
  .ZN(_2534_)
);

INV_X1 _6943_ (
  .A(_2534_),
  .ZN(_2535_)
);

NAND2_X2 _6944_ (
  .A1(_2501_),
  .A2(_2535_),
  .ZN(_2536_)
);

INV_X2 _6945_ (
  .A(_2536_),
  .ZN(_2537_)
);

NAND2_X1 _6946_ (
  .A1(_2466_),
  .A2(_2537_),
  .ZN(_2538_)
);

AND2_X2 _6947_ (
  .A1(_2537_),
  .A2(_2459_),
  .ZN(_2539_)
);

NAND2_X1 _6948_ (
  .A1(_2420_),
  .A2(_2539_),
  .ZN(_2540_)
);

NAND2_X1 _6949_ (
  .A1(_2504_),
  .A2(_2535_),
  .ZN(_2541_)
);

INV_X1 _6950_ (
  .A(_4355_),
  .ZN(_2542_)
);

OAI21_X1 _6951_ (
  .A(_2542_),
  .B1(_2528_),
  .B2(_2520_),
  .ZN(_2543_)
);

INV_X1 _6952_ (
  .A(_2543_),
  .ZN(_2544_)
);

NAND2_X1 _6953_ (
  .A1(_2541_),
  .A2(_2544_),
  .ZN(_2545_)
);

INV_X1 _6954_ (
  .A(_2545_),
  .ZN(_2546_)
);

NAND3_X2 _6955_ (
  .A1(_2538_),
  .A2(_2540_),
  .A3(_2546_),
  .ZN(_2547_)
);

INV_X1 _6956_ (
  .A(_2547_),
  .ZN(_2548_)
);

NOR2_X2 _6957_ (
  .A1(_0964_),
  .A2(\d_pipe[10][23] ),
  .ZN(_2549_)
);

NAND2_X4 _6958_ (
  .A1(_0949_),
  .A2(_2549_),
  .ZN(_2550_)
);

NAND2_X2 _6959_ (
  .A1(_2550_),
  .A2(_0638_),
  .ZN(_2551_)
);

INV_X1 _6960_ (
  .A(\s_pipe[10][23] ),
  .ZN(_2552_)
);

NAND2_X1 _6961_ (
  .A1(_2551_),
  .A2(_2552_),
  .ZN(_2553_)
);

NAND3_X1 _6962_ (
  .A1(_2550_),
  .A2(_0638_),
  .A3(\s_pipe[10][23] ),
  .ZN(_2554_)
);

NAND2_X1 _6963_ (
  .A1(_2553_),
  .A2(_2554_),
  .ZN(_2555_)
);

NAND2_X1 _6964_ (
  .A1(_2548_),
  .A2(_2555_),
  .ZN(_2556_)
);

NAND2_X1 _6965_ (
  .A1(_2551_),
  .A2(\s_pipe[10][23] ),
  .ZN(_2557_)
);

NAND3_X1 _6966_ (
  .A1(_2550_),
  .A2(_0638_),
  .A3(_2552_),
  .ZN(_2558_)
);

NAND2_X1 _6967_ (
  .A1(_2557_),
  .A2(_2558_),
  .ZN(_2559_)
);

NAND2_X1 _6968_ (
  .A1(_2559_),
  .A2(_2547_),
  .ZN(_2560_)
);

NAND3_X1 _6969_ (
  .A1(_2556_),
  .A2(_2560_),
  .A3(_2001_),
  .ZN(_2561_)
);

NAND2_X1 _6970_ (
  .A1(_1449_),
  .A2(\s_pipe[11][24] ),
  .ZN(_2562_)
);

NAND2_X1 _6971_ (
  .A1(_2561_),
  .A2(_2562_),
  .ZN(_0426_)
);

MUX2_X1 _6972_ (
  .A(\s_pipe[4][4] ),
  .B(\s_pipe[3][3] ),
  .S(_2066_),
  .Z(_0427_)
);

MUX2_X1 _6973_ (
  .A(\s_pipe[4][5] ),
  .B(\s_pipe[3][4] ),
  .S(_1565_),
  .Z(_0428_)
);

MUX2_X1 _6974_ (
  .A(\s_pipe[4][6] ),
  .B(\s_pipe[3][5] ),
  .S(_1566_),
  .Z(_0429_)
);

MUX2_X1 _6975_ (
  .A(\s_pipe[4][7] ),
  .B(\s_pipe[3][6] ),
  .S(_2068_),
  .Z(_0430_)
);

MUX2_X1 _6976_ (
  .A(\s_pipe[4][8] ),
  .B(\s_pipe[3][7] ),
  .S(_1861_),
  .Z(_0431_)
);

MUX2_X1 _6977_ (
  .A(\s_pipe[4][9] ),
  .B(\s_pipe[3][8] ),
  .S(_2007_),
  .Z(_0432_)
);

MUX2_X1 _6978_ (
  .A(\s_pipe[4][10] ),
  .B(\s_pipe[3][9] ),
  .S(_1933_),
  .Z(_0433_)
);

MUX2_X1 _6979_ (
  .A(\s_pipe[4][11] ),
  .B(\s_pipe[3][10] ),
  .S(_2067_),
  .Z(_0434_)
);

MUX2_X1 _6980_ (
  .A(\s_pipe[4][12] ),
  .B(_0125_),
  .S(_2068_),
  .Z(_0435_)
);

NAND2_X1 _6981_ (
  .A1(_1709_),
  .A2(\s_pipe[4][13] ),
  .ZN(_2563_)
);

OAI21_X1 _6982_ (
  .A(_2563_),
  .B1(_4053_),
  .B2(_1562_),
  .ZN(_0436_)
);

INV_X1 _6983_ (
  .A(_4052_),
  .ZN(_2564_)
);

NAND2_X1 _6984_ (
  .A1(_2564_),
  .A2(_4188_),
  .ZN(_2565_)
);

INV_X1 _6985_ (
  .A(_4188_),
  .ZN(_2566_)
);

NAND2_X1 _6986_ (
  .A1(_2566_),
  .A2(_4052_),
  .ZN(_2567_)
);

NAND3_X1 _6987_ (
  .A1(_2565_),
  .A2(_2567_),
  .A3(_1406_),
  .ZN(_2568_)
);

INV_X1 _6988_ (
  .A(\s_pipe[4][14] ),
  .ZN(_2569_)
);

OAI21_X1 _6989_ (
  .A(_2568_),
  .B1(_1408_),
  .B2(_2569_),
  .ZN(_0437_)
);

NOR2_X1 _6990_ (
  .A1(_2041_),
  .A2(\s_pipe[4][15] ),
  .ZN(_2570_)
);

INV_X1 _6991_ (
  .A(_4187_),
  .ZN(_2571_)
);

INV_X1 _6992_ (
  .A(_4184_),
  .ZN(_2572_)
);

OAI21_X2 _6993_ (
  .A(_2571_),
  .B1(_2566_),
  .B2(_2572_),
  .ZN(_2573_)
);

NAND2_X1 _6994_ (
  .A1(_4188_),
  .A2(_4185_),
  .ZN(_2574_)
);

NOR2_X1 _6995_ (
  .A1(_2574_),
  .A2(_4050_),
  .ZN(_2575_)
);

NOR2_X2 _6996_ (
  .A1(_2573_),
  .A2(_2575_),
  .ZN(_2576_)
);

INV_X1 _6997_ (
  .A(_4191_),
  .ZN(_2577_)
);

XNOR2_X1 _6998_ (
  .A(_2576_),
  .B(_2577_),
  .ZN(_2578_)
);

AOI21_X1 _6999_ (
  .A(_2570_),
  .B1(_2578_),
  .B2(_1363_),
  .ZN(_0438_)
);

NOR2_X1 _7000_ (
  .A1(_1364_),
  .A2(\s_pipe[4][16] ),
  .ZN(_2579_)
);

NOR2_X1 _7001_ (
  .A1(_4187_),
  .A2(_4190_),
  .ZN(_2580_)
);

INV_X1 _7002_ (
  .A(_4190_),
  .ZN(_2581_)
);

AOI22_X2 _7003_ (
  .A1(_2580_),
  .A2(_2565_),
  .B1(_2581_),
  .B2(_2577_),
  .ZN(_2582_)
);

BUF_X4 _7004_ (
  .A(_4194_),
  .Z(_2583_)
);

XNOR2_X1 _7005_ (
  .A(_2582_),
  .B(_2583_),
  .ZN(_2584_)
);

AOI21_X1 _7006_ (
  .A(_2579_),
  .B1(_2584_),
  .B2(_1363_),
  .ZN(_0439_)
);

NOR2_X1 _7007_ (
  .A1(_1353_),
  .A2(\s_pipe[4][17] ),
  .ZN(_2585_)
);

INV_X1 _7008_ (
  .A(_4193_),
  .ZN(_2586_)
);

INV_X1 _7009_ (
  .A(_2583_),
  .ZN(_2587_)
);

OAI21_X1 _7010_ (
  .A(_2586_),
  .B1(_2587_),
  .B2(_2581_),
  .ZN(_2588_)
);

INV_X1 _7011_ (
  .A(_2588_),
  .ZN(_2589_)
);

NAND2_X2 _7012_ (
  .A1(_4191_),
  .A2(_2583_),
  .ZN(_2590_)
);

OAI21_X1 _7013_ (
  .A(_2589_),
  .B1(_2576_),
  .B2(_2590_),
  .ZN(_2591_)
);

BUF_X4 _7014_ (
  .A(_4197_),
  .Z(_2592_)
);

XNOR2_X1 _7015_ (
  .A(_2591_),
  .B(_2592_),
  .ZN(_2593_)
);

AOI21_X1 _7016_ (
  .A(_2585_),
  .B1(_2593_),
  .B2(_1363_),
  .ZN(_0440_)
);

NOR2_X1 _7017_ (
  .A1(_2091_),
  .A2(\s_pipe[4][18] ),
  .ZN(_2594_)
);

INV_X1 _7018_ (
  .A(_4196_),
  .ZN(_2595_)
);

INV_X1 _7019_ (
  .A(_2592_),
  .ZN(_2596_)
);

OAI21_X2 _7020_ (
  .A(_2595_),
  .B1(_2596_),
  .B2(_2586_),
  .ZN(_2597_)
);

NAND2_X1 _7021_ (
  .A1(_2583_),
  .A2(_2592_),
  .ZN(_2598_)
);

INV_X1 _7022_ (
  .A(_2598_),
  .ZN(_2599_)
);

AOI21_X1 _7023_ (
  .A(_2597_),
  .B1(_2582_),
  .B2(_2599_),
  .ZN(_2600_)
);

INV_X1 _7024_ (
  .A(_4200_),
  .ZN(_2601_)
);

XNOR2_X1 _7025_ (
  .A(_2600_),
  .B(_2601_),
  .ZN(_2602_)
);

AOI21_X1 _7026_ (
  .A(_2594_),
  .B1(_2602_),
  .B2(_1381_),
  .ZN(_0441_)
);

INV_X1 _7027_ (
  .A(_2590_),
  .ZN(_2603_)
);

NAND2_X1 _7028_ (
  .A1(_2592_),
  .A2(_4200_),
  .ZN(_2604_)
);

INV_X1 _7029_ (
  .A(_2604_),
  .ZN(_2605_)
);

NAND2_X1 _7030_ (
  .A1(_2603_),
  .A2(_2605_),
  .ZN(_2606_)
);

OR2_X2 _7031_ (
  .A1(_2576_),
  .A2(_2606_),
  .ZN(_2607_)
);

NAND2_X1 _7032_ (
  .A1(_2588_),
  .A2(_2605_),
  .ZN(_2608_)
);

INV_X1 _7033_ (
  .A(_4199_),
  .ZN(_2609_)
);

OAI21_X1 _7034_ (
  .A(_2609_),
  .B1(_2601_),
  .B2(_2595_),
  .ZN(_2610_)
);

INV_X1 _7035_ (
  .A(_2610_),
  .ZN(_2611_)
);

NAND2_X1 _7036_ (
  .A1(_2608_),
  .A2(_2611_),
  .ZN(_2612_)
);

INV_X1 _7037_ (
  .A(_2612_),
  .ZN(_2613_)
);

NAND2_X1 _7038_ (
  .A1(_2607_),
  .A2(_2613_),
  .ZN(_2614_)
);

NAND2_X1 _7039_ (
  .A1(_2614_),
  .A2(_4203_),
  .ZN(_2615_)
);

INV_X1 _7040_ (
  .A(_4203_),
  .ZN(_2616_)
);

NAND3_X1 _7041_ (
  .A1(_2607_),
  .A2(_2613_),
  .A3(_2616_),
  .ZN(_2617_)
);

NAND3_X1 _7042_ (
  .A1(_2615_),
  .A2(_2617_),
  .A3(_1572_),
  .ZN(_2618_)
);

INV_X1 _7043_ (
  .A(\s_pipe[4][19] ),
  .ZN(_2619_)
);

OAI21_X1 _7044_ (
  .A(_2618_),
  .B1(_1408_),
  .B2(_2619_),
  .ZN(_0442_)
);

NAND2_X1 _7045_ (
  .A1(_4200_),
  .A2(_4203_),
  .ZN(_2620_)
);

NOR2_X2 _7046_ (
  .A1(_2598_),
  .A2(_2620_),
  .ZN(_2621_)
);

NAND2_X1 _7047_ (
  .A1(_2582_),
  .A2(_2621_),
  .ZN(_2622_)
);

INV_X1 _7048_ (
  .A(_2620_),
  .ZN(_2623_)
);

NAND2_X1 _7049_ (
  .A1(_2597_),
  .A2(_2623_),
  .ZN(_2624_)
);

INV_X1 _7050_ (
  .A(_4202_),
  .ZN(_2625_)
);

OAI21_X1 _7051_ (
  .A(_2625_),
  .B1(_2616_),
  .B2(_2609_),
  .ZN(_2626_)
);

INV_X1 _7052_ (
  .A(_2626_),
  .ZN(_2627_)
);

NAND2_X1 _7053_ (
  .A1(_2624_),
  .A2(_2627_),
  .ZN(_2628_)
);

INV_X1 _7054_ (
  .A(_2628_),
  .ZN(_2629_)
);

NAND2_X1 _7055_ (
  .A1(_2622_),
  .A2(_2629_),
  .ZN(_2630_)
);

NAND2_X1 _7056_ (
  .A1(_2630_),
  .A2(_4206_),
  .ZN(_2631_)
);

INV_X1 _7057_ (
  .A(_4206_),
  .ZN(_2632_)
);

NAND3_X1 _7058_ (
  .A1(_2622_),
  .A2(_2629_),
  .A3(_2632_),
  .ZN(_2633_)
);

NAND3_X1 _7059_ (
  .A1(_2631_),
  .A2(_2633_),
  .A3(_1572_),
  .ZN(_2634_)
);

INV_X1 _7060_ (
  .A(\s_pipe[4][20] ),
  .ZN(_2635_)
);

OAI21_X1 _7061_ (
  .A(_2634_),
  .B1(_1351_),
  .B2(_2635_),
  .ZN(_0443_)
);

NAND2_X1 _7062_ (
  .A1(_2573_),
  .A2(_2603_),
  .ZN(_2636_)
);

NAND2_X1 _7063_ (
  .A1(_2636_),
  .A2(_2589_),
  .ZN(_2637_)
);

NAND2_X1 _7064_ (
  .A1(_4203_),
  .A2(_4206_),
  .ZN(_2638_)
);

NOR2_X1 _7065_ (
  .A1(_2604_),
  .A2(_2638_),
  .ZN(_2639_)
);

NAND2_X1 _7066_ (
  .A1(_2637_),
  .A2(_2639_),
  .ZN(_2640_)
);

INV_X1 _7067_ (
  .A(_2638_),
  .ZN(_2641_)
);

NAND2_X1 _7068_ (
  .A1(_2610_),
  .A2(_2641_),
  .ZN(_2642_)
);

INV_X1 _7069_ (
  .A(_4205_),
  .ZN(_2643_)
);

OAI21_X1 _7070_ (
  .A(_2643_),
  .B1(_2632_),
  .B2(_2625_),
  .ZN(_2644_)
);

INV_X1 _7071_ (
  .A(_2644_),
  .ZN(_2645_)
);

NAND2_X1 _7072_ (
  .A1(_2642_),
  .A2(_2645_),
  .ZN(_2646_)
);

INV_X1 _7073_ (
  .A(_2646_),
  .ZN(_2647_)
);

NOR2_X1 _7074_ (
  .A1(_2574_),
  .A2(_2590_),
  .ZN(_2648_)
);

NAND3_X1 _7075_ (
  .A1(_2648_),
  .A2(_2639_),
  .A3(_4054_),
  .ZN(_2649_)
);

NAND3_X1 _7076_ (
  .A1(_2640_),
  .A2(_2647_),
  .A3(_2649_),
  .ZN(_2650_)
);

NAND2_X1 _7077_ (
  .A1(_2650_),
  .A2(_4209_),
  .ZN(_2651_)
);

INV_X1 _7078_ (
  .A(_4209_),
  .ZN(_2652_)
);

NAND4_X1 _7079_ (
  .A1(_2640_),
  .A2(_2649_),
  .A3(_2647_),
  .A4(_2652_),
  .ZN(_2653_)
);

NAND3_X1 _7080_ (
  .A1(_2651_),
  .A2(_2653_),
  .A3(_1669_),
  .ZN(_2654_)
);

NAND2_X1 _7081_ (
  .A1(_1449_),
  .A2(\s_pipe[4][21] ),
  .ZN(_2655_)
);

NAND2_X1 _7082_ (
  .A1(_2654_),
  .A2(_2655_),
  .ZN(_0444_)
);

OAI21_X1 _7083_ (
  .A(_2581_),
  .B1(_2577_),
  .B2(_2571_),
  .ZN(_2656_)
);

NAND2_X1 _7084_ (
  .A1(_2656_),
  .A2(_2599_),
  .ZN(_2657_)
);

INV_X1 _7085_ (
  .A(_2597_),
  .ZN(_2658_)
);

NAND2_X1 _7086_ (
  .A1(_2657_),
  .A2(_2658_),
  .ZN(_2659_)
);

NAND2_X1 _7087_ (
  .A1(_4206_),
  .A2(_4209_),
  .ZN(_2660_)
);

NOR2_X1 _7088_ (
  .A1(_2620_),
  .A2(_2660_),
  .ZN(_2661_)
);

NAND2_X1 _7089_ (
  .A1(_2659_),
  .A2(_2661_),
  .ZN(_2662_)
);

INV_X2 _7090_ (
  .A(_2660_),
  .ZN(_2663_)
);

NAND2_X1 _7091_ (
  .A1(_2626_),
  .A2(_2663_),
  .ZN(_2664_)
);

INV_X1 _7092_ (
  .A(_4208_),
  .ZN(_2665_)
);

OAI21_X1 _7093_ (
  .A(_2665_),
  .B1(_2652_),
  .B2(_2643_),
  .ZN(_2666_)
);

INV_X1 _7094_ (
  .A(_2666_),
  .ZN(_2667_)
);

NAND2_X1 _7095_ (
  .A1(_2664_),
  .A2(_2667_),
  .ZN(_2668_)
);

INV_X1 _7096_ (
  .A(_2668_),
  .ZN(_2669_)
);

NOR3_X1 _7097_ (
  .A1(_2598_),
  .A2(_2566_),
  .A3(_2577_),
  .ZN(_2670_)
);

NAND3_X1 _7098_ (
  .A1(_2670_),
  .A2(_2661_),
  .A3(_2564_),
  .ZN(_2671_)
);

NAND3_X1 _7099_ (
  .A1(_2662_),
  .A2(_2669_),
  .A3(_2671_),
  .ZN(_2672_)
);

NAND2_X1 _7100_ (
  .A1(_2672_),
  .A2(_4212_),
  .ZN(_2673_)
);

INV_X1 _7101_ (
  .A(_4212_),
  .ZN(_2674_)
);

NAND4_X1 _7102_ (
  .A1(_2662_),
  .A2(_2671_),
  .A3(_2669_),
  .A4(_2674_),
  .ZN(_2675_)
);

NAND3_X1 _7103_ (
  .A1(_2673_),
  .A2(_2675_),
  .A3(_2161_),
  .ZN(_2676_)
);

NAND2_X1 _7104_ (
  .A1(_1490_),
  .A2(\s_pipe[4][22] ),
  .ZN(_2677_)
);

NAND2_X1 _7105_ (
  .A1(_2676_),
  .A2(_2677_),
  .ZN(_0445_)
);

NAND2_X1 _7106_ (
  .A1(_4209_),
  .A2(_4212_),
  .ZN(_2678_)
);

OR2_X2 _7107_ (
  .A1(_2678_),
  .A2(_2638_),
  .ZN(_2679_)
);

INV_X1 _7108_ (
  .A(_2679_),
  .ZN(_2680_)
);

NAND2_X1 _7109_ (
  .A1(_2612_),
  .A2(_2680_),
  .ZN(_2681_)
);

INV_X1 _7110_ (
  .A(_4211_),
  .ZN(_2682_)
);

OAI21_X1 _7111_ (
  .A(_2682_),
  .B1(_2674_),
  .B2(_2665_),
  .ZN(_2683_)
);

INV_X1 _7112_ (
  .A(_2683_),
  .ZN(_2684_)
);

OAI21_X1 _7113_ (
  .A(_2684_),
  .B1(_2645_),
  .B2(_2678_),
  .ZN(_2685_)
);

INV_X1 _7114_ (
  .A(_2685_),
  .ZN(_2686_)
);

INV_X1 _7115_ (
  .A(_2576_),
  .ZN(_2687_)
);

NOR2_X2 _7116_ (
  .A1(_2679_),
  .A2(_2606_),
  .ZN(_2688_)
);

NAND2_X1 _7117_ (
  .A1(_2687_),
  .A2(_2688_),
  .ZN(_2689_)
);

INV_X1 _7118_ (
  .A(_4215_),
  .ZN(_2690_)
);

NAND4_X1 _7119_ (
  .A1(_2681_),
  .A2(_2686_),
  .A3(_2689_),
  .A4(_2690_),
  .ZN(_2691_)
);

NAND3_X1 _7120_ (
  .A1(_2681_),
  .A2(_2686_),
  .A3(_2689_),
  .ZN(_2692_)
);

NAND2_X1 _7121_ (
  .A1(_2692_),
  .A2(_4215_),
  .ZN(_2693_)
);

NAND3_X1 _7122_ (
  .A1(_2691_),
  .A2(_2693_),
  .A3(_1669_),
  .ZN(_2694_)
);

NAND2_X1 _7123_ (
  .A1(_1490_),
  .A2(\s_pipe[4][23] ),
  .ZN(_2695_)
);

NAND2_X1 _7124_ (
  .A1(_2694_),
  .A2(_2695_),
  .ZN(_0446_)
);

NAND2_X1 _7125_ (
  .A1(_4212_),
  .A2(_4215_),
  .ZN(_2696_)
);

INV_X1 _7126_ (
  .A(_2696_),
  .ZN(_2697_)
);

NAND2_X1 _7127_ (
  .A1(_2663_),
  .A2(_2697_),
  .ZN(_2698_)
);

INV_X2 _7128_ (
  .A(_2698_),
  .ZN(_2699_)
);

NAND2_X1 _7129_ (
  .A1(_2628_),
  .A2(_2699_),
  .ZN(_2700_)
);

AND2_X2 _7130_ (
  .A1(_2699_),
  .A2(_2621_),
  .ZN(_2701_)
);

NAND2_X2 _7131_ (
  .A1(_2582_),
  .A2(_2701_),
  .ZN(_2702_)
);

NAND2_X1 _7132_ (
  .A1(_2666_),
  .A2(_2697_),
  .ZN(_2703_)
);

INV_X1 _7133_ (
  .A(_4214_),
  .ZN(_2704_)
);

OAI21_X1 _7134_ (
  .A(_2704_),
  .B1(_2690_),
  .B2(_2682_),
  .ZN(_2705_)
);

INV_X1 _7135_ (
  .A(_2705_),
  .ZN(_2706_)
);

NAND2_X1 _7136_ (
  .A1(_2703_),
  .A2(_2706_),
  .ZN(_2707_)
);

INV_X1 _7137_ (
  .A(_2707_),
  .ZN(_2708_)
);

NAND3_X2 _7138_ (
  .A1(_2700_),
  .A2(_2702_),
  .A3(_2708_),
  .ZN(_2709_)
);

INV_X1 _7139_ (
  .A(_2709_),
  .ZN(_2710_)
);

NOR2_X2 _7140_ (
  .A1(_0795_),
  .A2(\d_pipe[3][23] ),
  .ZN(_2711_)
);

NAND2_X4 _7141_ (
  .A1(_0779_),
  .A2(_2711_),
  .ZN(_2712_)
);

NAND2_X2 _7142_ (
  .A1(_2712_),
  .A2(_0629_),
  .ZN(_2713_)
);

INV_X1 _7143_ (
  .A(\s_pipe[3][23] ),
  .ZN(_2714_)
);

NAND2_X1 _7144_ (
  .A1(_2713_),
  .A2(_2714_),
  .ZN(_2715_)
);

NAND3_X1 _7145_ (
  .A1(_2712_),
  .A2(_0629_),
  .A3(\s_pipe[3][23] ),
  .ZN(_2716_)
);

NAND2_X1 _7146_ (
  .A1(_2715_),
  .A2(_2716_),
  .ZN(_2717_)
);

NAND2_X1 _7147_ (
  .A1(_2710_),
  .A2(_2717_),
  .ZN(_2718_)
);

NAND2_X1 _7148_ (
  .A1(_2713_),
  .A2(\s_pipe[3][23] ),
  .ZN(_2719_)
);

NAND3_X1 _7149_ (
  .A1(_2712_),
  .A2(_0629_),
  .A3(_2714_),
  .ZN(_2720_)
);

NAND2_X1 _7150_ (
  .A1(_2719_),
  .A2(_2720_),
  .ZN(_2721_)
);

NAND2_X1 _7151_ (
  .A1(_2721_),
  .A2(_2709_),
  .ZN(_2722_)
);

NAND3_X1 _7152_ (
  .A1(_2718_),
  .A2(_2722_),
  .A3(_2349_),
  .ZN(_2723_)
);

NAND2_X1 _7153_ (
  .A1(_1490_),
  .A2(\s_pipe[4][24] ),
  .ZN(_2724_)
);

NAND2_X1 _7154_ (
  .A1(_2723_),
  .A2(_2724_),
  .ZN(_0447_)
);

NAND2_X1 _7155_ (
  .A1(_2057_),
  .A2(\s_pipe[9][9] ),
  .ZN(_2725_)
);

INV_X1 _7156_ (
  .A(\s_pipe[8][8] ),
  .ZN(_2726_)
);

OAI21_X1 _7157_ (
  .A(_2725_),
  .B1(_1524_),
  .B2(_2726_),
  .ZN(_0448_)
);

NAND2_X1 _7158_ (
  .A1(_2057_),
  .A2(\s_pipe[9][10] ),
  .ZN(_2727_)
);

INV_X1 _7159_ (
  .A(\s_pipe[8][9] ),
  .ZN(_2728_)
);

OAI21_X1 _7160_ (
  .A(_2727_),
  .B1(_1865_),
  .B2(_2728_),
  .ZN(_0449_)
);

NAND2_X1 _7161_ (
  .A1(_2057_),
  .A2(\s_pipe[9][11] ),
  .ZN(_2729_)
);

INV_X1 _7162_ (
  .A(\s_pipe[8][10] ),
  .ZN(_2730_)
);

OAI21_X1 _7163_ (
  .A(_2729_),
  .B1(_1524_),
  .B2(_2730_),
  .ZN(_0450_)
);

MUX2_X1 _7164_ (
  .A(\s_pipe[9][12] ),
  .B(_0130_),
  .S(_1934_),
  .Z(_0451_)
);

NAND2_X1 _7165_ (
  .A1(_2057_),
  .A2(\s_pipe[9][13] ),
  .ZN(_2731_)
);

OAI21_X1 _7166_ (
  .A(_2731_),
  .B1(_4091_),
  .B2(_2054_),
  .ZN(_0452_)
);

INV_X1 _7167_ (
  .A(_4090_),
  .ZN(_2732_)
);

NAND2_X1 _7168_ (
  .A1(_2732_),
  .A2(_4401_),
  .ZN(_2733_)
);

INV_X1 _7169_ (
  .A(_4401_),
  .ZN(_2734_)
);

NAND2_X1 _7170_ (
  .A1(_2734_),
  .A2(_4090_),
  .ZN(_2735_)
);

NAND3_X1 _7171_ (
  .A1(_2733_),
  .A2(_2735_),
  .A3(_2238_),
  .ZN(_2736_)
);

INV_X1 _7172_ (
  .A(\s_pipe[9][14] ),
  .ZN(_2737_)
);

OAI21_X1 _7173_ (
  .A(_2736_),
  .B1(_2291_),
  .B2(_2737_),
  .ZN(_0453_)
);

NOR2_X1 _7174_ (
  .A1(_1364_),
  .A2(_0134_),
  .ZN(_2738_)
);

INV_X1 _7175_ (
  .A(_4400_),
  .ZN(_2739_)
);

INV_X1 _7176_ (
  .A(_4397_),
  .ZN(_2740_)
);

OAI21_X2 _7177_ (
  .A(_2739_),
  .B1(_2734_),
  .B2(_2740_),
  .ZN(_2741_)
);

NAND2_X1 _7178_ (
  .A1(_4401_),
  .A2(_4398_),
  .ZN(_2742_)
);

NOR2_X1 _7179_ (
  .A1(_2742_),
  .A2(_4089_),
  .ZN(_2743_)
);

NOR2_X2 _7180_ (
  .A1(_2741_),
  .A2(_2743_),
  .ZN(_2744_)
);

INV_X1 _7181_ (
  .A(_4404_),
  .ZN(_2745_)
);

XNOR2_X1 _7182_ (
  .A(_2744_),
  .B(_2745_),
  .ZN(_2746_)
);

AOI21_X1 _7183_ (
  .A(_2738_),
  .B1(_2746_),
  .B2(_1587_),
  .ZN(_0454_)
);

NOR2_X1 _7184_ (
  .A1(_1353_),
  .A2(_0135_),
  .ZN(_2747_)
);

NOR2_X1 _7185_ (
  .A1(_4400_),
  .A2(_4403_),
  .ZN(_2748_)
);

INV_X1 _7186_ (
  .A(_4403_),
  .ZN(_2749_)
);

AOI22_X2 _7187_ (
  .A1(_2748_),
  .A2(_2733_),
  .B1(_2749_),
  .B2(_2745_),
  .ZN(_2750_)
);

BUF_X4 _7188_ (
  .A(_4407_),
  .Z(_2751_)
);

XNOR2_X1 _7189_ (
  .A(_2750_),
  .B(_2751_),
  .ZN(_2752_)
);

AOI21_X1 _7190_ (
  .A(_2747_),
  .B1(_2752_),
  .B2(_2265_),
  .ZN(_0455_)
);

NOR2_X1 _7191_ (
  .A1(_2041_),
  .A2(_0136_),
  .ZN(_2753_)
);

INV_X1 _7192_ (
  .A(_4406_),
  .ZN(_2754_)
);

INV_X1 _7193_ (
  .A(_2751_),
  .ZN(_2755_)
);

OAI21_X1 _7194_ (
  .A(_2754_),
  .B1(_2755_),
  .B2(_2749_),
  .ZN(_2756_)
);

INV_X1 _7195_ (
  .A(_2756_),
  .ZN(_2757_)
);

NAND2_X2 _7196_ (
  .A1(_4404_),
  .A2(_2751_),
  .ZN(_2758_)
);

OAI21_X1 _7197_ (
  .A(_2757_),
  .B1(_2744_),
  .B2(_2758_),
  .ZN(_2759_)
);

BUF_X4 _7198_ (
  .A(_4410_),
  .Z(_2760_)
);

XNOR2_X1 _7199_ (
  .A(_2759_),
  .B(_2760_),
  .ZN(_2761_)
);

AOI21_X1 _7200_ (
  .A(_2753_),
  .B1(_2761_),
  .B2(_2265_),
  .ZN(_0456_)
);

NOR2_X1 _7201_ (
  .A1(_2041_),
  .A2(_0137_),
  .ZN(_2762_)
);

INV_X1 _7202_ (
  .A(_4409_),
  .ZN(_2763_)
);

INV_X1 _7203_ (
  .A(_2760_),
  .ZN(_2764_)
);

OAI21_X2 _7204_ (
  .A(_2763_),
  .B1(_2764_),
  .B2(_2754_),
  .ZN(_2765_)
);

NAND2_X1 _7205_ (
  .A1(_2751_),
  .A2(_2760_),
  .ZN(_2766_)
);

INV_X1 _7206_ (
  .A(_2766_),
  .ZN(_2767_)
);

AOI21_X1 _7207_ (
  .A(_2765_),
  .B1(_2750_),
  .B2(_2767_),
  .ZN(_2768_)
);

INV_X1 _7208_ (
  .A(_4413_),
  .ZN(_2769_)
);

XNOR2_X1 _7209_ (
  .A(_2768_),
  .B(_2769_),
  .ZN(_2770_)
);

AOI21_X1 _7210_ (
  .A(_2762_),
  .B1(_2770_),
  .B2(_2265_),
  .ZN(_0457_)
);

INV_X1 _7211_ (
  .A(_2758_),
  .ZN(_2771_)
);

NAND2_X1 _7212_ (
  .A1(_2760_),
  .A2(_4413_),
  .ZN(_2772_)
);

INV_X1 _7213_ (
  .A(_2772_),
  .ZN(_2773_)
);

NAND2_X1 _7214_ (
  .A1(_2771_),
  .A2(_2773_),
  .ZN(_2774_)
);

OR2_X2 _7215_ (
  .A1(_2744_),
  .A2(_2774_),
  .ZN(_2775_)
);

NAND2_X1 _7216_ (
  .A1(_2756_),
  .A2(_2773_),
  .ZN(_2776_)
);

INV_X1 _7217_ (
  .A(_4412_),
  .ZN(_2777_)
);

OAI21_X1 _7218_ (
  .A(_2777_),
  .B1(_2769_),
  .B2(_2763_),
  .ZN(_2778_)
);

INV_X1 _7219_ (
  .A(_2778_),
  .ZN(_2779_)
);

NAND2_X1 _7220_ (
  .A1(_2776_),
  .A2(_2779_),
  .ZN(_2780_)
);

INV_X1 _7221_ (
  .A(_2780_),
  .ZN(_2781_)
);

NAND2_X1 _7222_ (
  .A1(_2775_),
  .A2(_2781_),
  .ZN(_2782_)
);

NAND2_X1 _7223_ (
  .A1(_2782_),
  .A2(_4416_),
  .ZN(_2783_)
);

INV_X1 _7224_ (
  .A(_4416_),
  .ZN(_2784_)
);

NAND3_X1 _7225_ (
  .A1(_2775_),
  .A2(_2781_),
  .A3(_2784_),
  .ZN(_2785_)
);

NAND3_X1 _7226_ (
  .A1(_2783_),
  .A2(_2785_),
  .A3(_1348_),
  .ZN(_2786_)
);

INV_X1 _7227_ (
  .A(_0138_),
  .ZN(_2787_)
);

OAI21_X1 _7228_ (
  .A(_2786_),
  .B1(_1901_),
  .B2(_2787_),
  .ZN(_0458_)
);

NAND2_X1 _7229_ (
  .A1(_4413_),
  .A2(_4416_),
  .ZN(_2788_)
);

NOR2_X2 _7230_ (
  .A1(_2766_),
  .A2(_2788_),
  .ZN(_2789_)
);

NAND2_X1 _7231_ (
  .A1(_2750_),
  .A2(_2789_),
  .ZN(_2790_)
);

INV_X1 _7232_ (
  .A(_2788_),
  .ZN(_2791_)
);

NAND2_X1 _7233_ (
  .A1(_2765_),
  .A2(_2791_),
  .ZN(_2792_)
);

INV_X1 _7234_ (
  .A(_4415_),
  .ZN(_2793_)
);

OAI21_X1 _7235_ (
  .A(_2793_),
  .B1(_2784_),
  .B2(_2777_),
  .ZN(_2794_)
);

INV_X1 _7236_ (
  .A(_2794_),
  .ZN(_2795_)
);

NAND2_X1 _7237_ (
  .A1(_2792_),
  .A2(_2795_),
  .ZN(_2796_)
);

INV_X1 _7238_ (
  .A(_2796_),
  .ZN(_2797_)
);

NAND2_X1 _7239_ (
  .A1(_2790_),
  .A2(_2797_),
  .ZN(_2798_)
);

NAND2_X1 _7240_ (
  .A1(_2798_),
  .A2(_4419_),
  .ZN(_2799_)
);

INV_X1 _7241_ (
  .A(_4419_),
  .ZN(_2800_)
);

NAND3_X1 _7242_ (
  .A1(_2790_),
  .A2(_2797_),
  .A3(_2800_),
  .ZN(_2801_)
);

NAND3_X1 _7243_ (
  .A1(_2799_),
  .A2(_2801_),
  .A3(_1572_),
  .ZN(_2802_)
);

INV_X1 _7244_ (
  .A(_0139_),
  .ZN(_2803_)
);

OAI21_X1 _7245_ (
  .A(_2802_),
  .B1(_1351_),
  .B2(_2803_),
  .ZN(_0459_)
);

NAND2_X1 _7246_ (
  .A1(_2741_),
  .A2(_2771_),
  .ZN(_2804_)
);

NAND2_X1 _7247_ (
  .A1(_2804_),
  .A2(_2757_),
  .ZN(_2805_)
);

NAND2_X1 _7248_ (
  .A1(_4416_),
  .A2(_4419_),
  .ZN(_2806_)
);

NOR2_X1 _7249_ (
  .A1(_2772_),
  .A2(_2806_),
  .ZN(_2807_)
);

NAND2_X1 _7250_ (
  .A1(_2805_),
  .A2(_2807_),
  .ZN(_2808_)
);

INV_X1 _7251_ (
  .A(_2806_),
  .ZN(_2809_)
);

NAND2_X1 _7252_ (
  .A1(_2778_),
  .A2(_2809_),
  .ZN(_2810_)
);

INV_X1 _7253_ (
  .A(_4418_),
  .ZN(_2811_)
);

OAI21_X1 _7254_ (
  .A(_2811_),
  .B1(_2800_),
  .B2(_2793_),
  .ZN(_2812_)
);

INV_X1 _7255_ (
  .A(_2812_),
  .ZN(_2813_)
);

NAND2_X1 _7256_ (
  .A1(_2810_),
  .A2(_2813_),
  .ZN(_2814_)
);

INV_X1 _7257_ (
  .A(_2814_),
  .ZN(_2815_)
);

NOR2_X1 _7258_ (
  .A1(_2742_),
  .A2(_2758_),
  .ZN(_2816_)
);

NAND3_X1 _7259_ (
  .A1(_2816_),
  .A2(_2807_),
  .A3(_4093_),
  .ZN(_2817_)
);

NAND3_X1 _7260_ (
  .A1(_2808_),
  .A2(_2815_),
  .A3(_2817_),
  .ZN(_2818_)
);

NAND2_X1 _7261_ (
  .A1(_2818_),
  .A2(_4422_),
  .ZN(_2819_)
);

INV_X1 _7262_ (
  .A(_4422_),
  .ZN(_2820_)
);

NAND4_X1 _7263_ (
  .A1(_2808_),
  .A2(_2817_),
  .A3(_2815_),
  .A4(_2820_),
  .ZN(_2821_)
);

NAND3_X1 _7264_ (
  .A1(_2819_),
  .A2(_2821_),
  .A3(_2349_),
  .ZN(_2822_)
);

NAND2_X1 _7265_ (
  .A1(_1728_),
  .A2(_0131_),
  .ZN(_2823_)
);

NAND2_X1 _7266_ (
  .A1(_2822_),
  .A2(_2823_),
  .ZN(_0460_)
);

OAI21_X1 _7267_ (
  .A(_2749_),
  .B1(_2745_),
  .B2(_2739_),
  .ZN(_2824_)
);

NAND2_X1 _7268_ (
  .A1(_2824_),
  .A2(_2767_),
  .ZN(_2825_)
);

INV_X1 _7269_ (
  .A(_2765_),
  .ZN(_2826_)
);

NAND2_X1 _7270_ (
  .A1(_2825_),
  .A2(_2826_),
  .ZN(_2827_)
);

NAND2_X2 _7271_ (
  .A1(_4419_),
  .A2(_4422_),
  .ZN(_2828_)
);

NOR2_X1 _7272_ (
  .A1(_2788_),
  .A2(_2828_),
  .ZN(_2829_)
);

NAND2_X1 _7273_ (
  .A1(_2827_),
  .A2(_2829_),
  .ZN(_2830_)
);

INV_X2 _7274_ (
  .A(_2828_),
  .ZN(_2831_)
);

NAND2_X1 _7275_ (
  .A1(_2794_),
  .A2(_2831_),
  .ZN(_2832_)
);

INV_X1 _7276_ (
  .A(_4421_),
  .ZN(_2833_)
);

OAI21_X1 _7277_ (
  .A(_2833_),
  .B1(_2820_),
  .B2(_2811_),
  .ZN(_2834_)
);

INV_X1 _7278_ (
  .A(_2834_),
  .ZN(_2835_)
);

NAND2_X1 _7279_ (
  .A1(_2832_),
  .A2(_2835_),
  .ZN(_2836_)
);

INV_X1 _7280_ (
  .A(_2836_),
  .ZN(_2837_)
);

NOR3_X1 _7281_ (
  .A1(_2766_),
  .A2(_2734_),
  .A3(_2745_),
  .ZN(_2838_)
);

NAND3_X1 _7282_ (
  .A1(_2838_),
  .A2(_2829_),
  .A3(_2732_),
  .ZN(_2839_)
);

NAND3_X1 _7283_ (
  .A1(_2830_),
  .A2(_2837_),
  .A3(_2839_),
  .ZN(_2840_)
);

NAND2_X1 _7284_ (
  .A1(_2840_),
  .A2(_4425_),
  .ZN(_2841_)
);

INV_X1 _7285_ (
  .A(_4425_),
  .ZN(_2842_)
);

NAND4_X1 _7286_ (
  .A1(_2830_),
  .A2(_2839_),
  .A3(_2837_),
  .A4(_2842_),
  .ZN(_2843_)
);

NAND3_X1 _7287_ (
  .A1(_2841_),
  .A2(_2843_),
  .A3(_2161_),
  .ZN(_2844_)
);

NAND2_X1 _7288_ (
  .A1(_1859_),
  .A2(_0132_),
  .ZN(_2845_)
);

NAND2_X1 _7289_ (
  .A1(_2844_),
  .A2(_2845_),
  .ZN(_0461_)
);

NAND2_X1 _7290_ (
  .A1(_4422_),
  .A2(_4425_),
  .ZN(_2846_)
);

OR2_X2 _7291_ (
  .A1(_2846_),
  .A2(_2806_),
  .ZN(_2847_)
);

INV_X1 _7292_ (
  .A(_2847_),
  .ZN(_2848_)
);

NAND2_X1 _7293_ (
  .A1(_2780_),
  .A2(_2848_),
  .ZN(_2849_)
);

INV_X1 _7294_ (
  .A(_4424_),
  .ZN(_2850_)
);

OAI21_X1 _7295_ (
  .A(_2850_),
  .B1(_2842_),
  .B2(_2833_),
  .ZN(_2851_)
);

INV_X1 _7296_ (
  .A(_2851_),
  .ZN(_2852_)
);

OAI21_X1 _7297_ (
  .A(_2852_),
  .B1(_2813_),
  .B2(_2846_),
  .ZN(_2853_)
);

INV_X1 _7298_ (
  .A(_2853_),
  .ZN(_2854_)
);

INV_X1 _7299_ (
  .A(_2744_),
  .ZN(_2855_)
);

NOR2_X2 _7300_ (
  .A1(_2847_),
  .A2(_2774_),
  .ZN(_2856_)
);

NAND2_X1 _7301_ (
  .A1(_2855_),
  .A2(_2856_),
  .ZN(_2857_)
);

INV_X1 _7302_ (
  .A(_4428_),
  .ZN(_2858_)
);

NAND4_X1 _7303_ (
  .A1(_2849_),
  .A2(_2854_),
  .A3(_2857_),
  .A4(_2858_),
  .ZN(_2859_)
);

NAND3_X1 _7304_ (
  .A1(_2849_),
  .A2(_2854_),
  .A3(_2857_),
  .ZN(_2860_)
);

NAND2_X1 _7305_ (
  .A1(_2860_),
  .A2(_4428_),
  .ZN(_2861_)
);

NAND3_X1 _7306_ (
  .A1(_2859_),
  .A2(_2861_),
  .A3(_2161_),
  .ZN(_2862_)
);

NAND2_X1 _7307_ (
  .A1(_1859_),
  .A2(_0133_),
  .ZN(_2863_)
);

NAND2_X1 _7308_ (
  .A1(_2862_),
  .A2(_2863_),
  .ZN(_0462_)
);

NAND2_X1 _7309_ (
  .A1(_4425_),
  .A2(_4428_),
  .ZN(_2864_)
);

INV_X1 _7310_ (
  .A(_2864_),
  .ZN(_2865_)
);

NAND2_X1 _7311_ (
  .A1(_2831_),
  .A2(_2865_),
  .ZN(_2866_)
);

INV_X2 _7312_ (
  .A(_2866_),
  .ZN(_2867_)
);

NAND2_X1 _7313_ (
  .A1(_2796_),
  .A2(_2867_),
  .ZN(_2868_)
);

AND2_X2 _7314_ (
  .A1(_2867_),
  .A2(_2789_),
  .ZN(_2869_)
);

NAND2_X1 _7315_ (
  .A1(_2750_),
  .A2(_2869_),
  .ZN(_2870_)
);

NAND2_X1 _7316_ (
  .A1(_2834_),
  .A2(_2865_),
  .ZN(_2871_)
);

INV_X1 _7317_ (
  .A(_4427_),
  .ZN(_2872_)
);

OAI21_X1 _7318_ (
  .A(_2872_),
  .B1(_2858_),
  .B2(_2850_),
  .ZN(_2873_)
);

INV_X1 _7319_ (
  .A(_2873_),
  .ZN(_2874_)
);

NAND2_X1 _7320_ (
  .A1(_2871_),
  .A2(_2874_),
  .ZN(_2875_)
);

INV_X1 _7321_ (
  .A(_2875_),
  .ZN(_2876_)
);

NAND3_X2 _7322_ (
  .A1(_2868_),
  .A2(_2870_),
  .A3(_2876_),
  .ZN(_2877_)
);

INV_X1 _7323_ (
  .A(_2877_),
  .ZN(_2878_)
);

NOR2_X2 _7324_ (
  .A1(_1077_),
  .A2(\d_pipe[8][23] ),
  .ZN(_2879_)
);

NAND2_X4 _7325_ (
  .A1(_1061_),
  .A2(_2879_),
  .ZN(_2880_)
);

NAND2_X2 _7326_ (
  .A1(_2880_),
  .A2(_0645_),
  .ZN(_2881_)
);

INV_X1 _7327_ (
  .A(\s_pipe[8][23] ),
  .ZN(_2882_)
);

NAND2_X1 _7328_ (
  .A1(_2881_),
  .A2(_2882_),
  .ZN(_2883_)
);

NAND3_X1 _7329_ (
  .A1(_2880_),
  .A2(_0645_),
  .A3(\s_pipe[8][23] ),
  .ZN(_2884_)
);

NAND2_X1 _7330_ (
  .A1(_2883_),
  .A2(_2884_),
  .ZN(_2885_)
);

NAND2_X1 _7331_ (
  .A1(_2878_),
  .A2(_2885_),
  .ZN(_2886_)
);

NAND2_X1 _7332_ (
  .A1(_2881_),
  .A2(\s_pipe[8][23] ),
  .ZN(_2887_)
);

NAND3_X1 _7333_ (
  .A1(_2880_),
  .A2(_0645_),
  .A3(_2882_),
  .ZN(_2888_)
);

NAND2_X1 _7334_ (
  .A1(_2887_),
  .A2(_2888_),
  .ZN(_2889_)
);

NAND2_X1 _7335_ (
  .A1(_2889_),
  .A2(_2877_),
  .ZN(_2890_)
);

NAND3_X1 _7336_ (
  .A1(_2886_),
  .A2(_2890_),
  .A3(_2161_),
  .ZN(_2891_)
);

NAND2_X1 _7337_ (
  .A1(_1859_),
  .A2(_0641_),
  .ZN(_2892_)
);

NAND2_X1 _7338_ (
  .A1(_2891_),
  .A2(_2892_),
  .ZN(_0463_)
);

MUX2_X1 _7339_ (
  .A(\s_pipe[5][5] ),
  .B(\s_pipe[4][4] ),
  .S(_2066_),
  .Z(_0464_)
);

MUX2_X1 _7340_ (
  .A(\s_pipe[5][6] ),
  .B(\s_pipe[4][5] ),
  .S(_2007_),
  .Z(_0465_)
);

MUX2_X1 _7341_ (
  .A(\s_pipe[5][7] ),
  .B(\s_pipe[4][6] ),
  .S(_1565_),
  .Z(_0466_)
);

MUX2_X1 _7342_ (
  .A(\s_pipe[5][8] ),
  .B(\s_pipe[4][7] ),
  .S(_2007_),
  .Z(_0467_)
);

MUX2_X1 _7343_ (
  .A(\s_pipe[5][9] ),
  .B(\s_pipe[4][8] ),
  .S(_2041_),
  .Z(_0468_)
);

MUX2_X1 _7344_ (
  .A(\s_pipe[5][10] ),
  .B(\s_pipe[4][9] ),
  .S(_2041_),
  .Z(_0469_)
);

MUX2_X1 _7345_ (
  .A(\s_pipe[5][11] ),
  .B(\s_pipe[4][10] ),
  .S(_1952_),
  .Z(_0470_)
);

MUX2_X1 _7346_ (
  .A(\s_pipe[5][12] ),
  .B(_0126_),
  .S(_2041_),
  .Z(_0471_)
);

NAND2_X1 _7347_ (
  .A1(_1881_),
  .A2(\s_pipe[5][13] ),
  .ZN(_2893_)
);

OAI21_X1 _7348_ (
  .A(_2893_),
  .B1(_4119_),
  .B2(_2054_),
  .ZN(_0472_)
);

INV_X1 _7349_ (
  .A(_4118_),
  .ZN(_2894_)
);

NAND2_X1 _7350_ (
  .A1(_2894_),
  .A2(_4545_),
  .ZN(_2895_)
);

INV_X1 _7351_ (
  .A(_4545_),
  .ZN(_2896_)
);

NAND2_X1 _7352_ (
  .A1(_2896_),
  .A2(_4118_),
  .ZN(_2897_)
);

NAND3_X1 _7353_ (
  .A1(_2895_),
  .A2(_2897_),
  .A3(_1348_),
  .ZN(_2898_)
);

INV_X1 _7354_ (
  .A(\s_pipe[5][14] ),
  .ZN(_2899_)
);

OAI21_X1 _7355_ (
  .A(_2898_),
  .B1(_1548_),
  .B2(_2899_),
  .ZN(_0473_)
);

NOR2_X1 _7356_ (
  .A1(_1371_),
  .A2(\s_pipe[5][15] ),
  .ZN(_2900_)
);

INV_X1 _7357_ (
  .A(_4544_),
  .ZN(_2901_)
);

INV_X1 _7358_ (
  .A(_4541_),
  .ZN(_2902_)
);

OAI21_X2 _7359_ (
  .A(_2901_),
  .B1(_2896_),
  .B2(_2902_),
  .ZN(_2903_)
);

NAND2_X1 _7360_ (
  .A1(_4545_),
  .A2(_4542_),
  .ZN(_2904_)
);

NOR2_X1 _7361_ (
  .A1(_2904_),
  .A2(_4117_),
  .ZN(_2905_)
);

NOR2_X2 _7362_ (
  .A1(_2903_),
  .A2(_2905_),
  .ZN(_2906_)
);

INV_X1 _7363_ (
  .A(_4548_),
  .ZN(_2907_)
);

XNOR2_X1 _7364_ (
  .A(_2906_),
  .B(_2907_),
  .ZN(_2908_)
);

AOI21_X1 _7365_ (
  .A(_2900_),
  .B1(_2908_),
  .B2(_2265_),
  .ZN(_0474_)
);

NOR2_X1 _7366_ (
  .A1(_1353_),
  .A2(\s_pipe[5][16] ),
  .ZN(_2909_)
);

NOR2_X1 _7367_ (
  .A1(_4544_),
  .A2(_4547_),
  .ZN(_2910_)
);

INV_X1 _7368_ (
  .A(_4547_),
  .ZN(_2911_)
);

AOI22_X2 _7369_ (
  .A1(_2910_),
  .A2(_2895_),
  .B1(_2911_),
  .B2(_2907_),
  .ZN(_2912_)
);

BUF_X4 _7370_ (
  .A(_4551_),
  .Z(_2913_)
);

XNOR2_X1 _7371_ (
  .A(_2912_),
  .B(_2913_),
  .ZN(_2914_)
);

AOI21_X1 _7372_ (
  .A(_2909_),
  .B1(_2914_),
  .B2(_2265_),
  .ZN(_0475_)
);

NOR2_X1 _7373_ (
  .A1(_2041_),
  .A2(\s_pipe[5][17] ),
  .ZN(_2915_)
);

INV_X1 _7374_ (
  .A(_4550_),
  .ZN(_2916_)
);

INV_X1 _7375_ (
  .A(_2913_),
  .ZN(_2917_)
);

OAI21_X1 _7376_ (
  .A(_2916_),
  .B1(_2917_),
  .B2(_2911_),
  .ZN(_2918_)
);

INV_X1 _7377_ (
  .A(_2918_),
  .ZN(_2919_)
);

NAND2_X2 _7378_ (
  .A1(_4548_),
  .A2(_2913_),
  .ZN(_2920_)
);

OAI21_X1 _7379_ (
  .A(_2919_),
  .B1(_2906_),
  .B2(_2920_),
  .ZN(_2921_)
);

BUF_X2 _7380_ (
  .A(_4554_),
  .Z(_2922_)
);

XNOR2_X1 _7381_ (
  .A(_2921_),
  .B(_2922_),
  .ZN(_2923_)
);

AOI21_X1 _7382_ (
  .A(_2915_),
  .B1(_2923_),
  .B2(_2265_),
  .ZN(_0476_)
);

NOR2_X1 _7383_ (
  .A1(_2041_),
  .A2(\s_pipe[5][18] ),
  .ZN(_2924_)
);

INV_X1 _7384_ (
  .A(_4553_),
  .ZN(_2925_)
);

INV_X1 _7385_ (
  .A(_2922_),
  .ZN(_2926_)
);

OAI21_X2 _7386_ (
  .A(_2925_),
  .B1(_2926_),
  .B2(_2916_),
  .ZN(_2927_)
);

NAND2_X1 _7387_ (
  .A1(_2913_),
  .A2(_2922_),
  .ZN(_2928_)
);

INV_X1 _7388_ (
  .A(_2928_),
  .ZN(_2929_)
);

AOI21_X1 _7389_ (
  .A(_2927_),
  .B1(_2912_),
  .B2(_2929_),
  .ZN(_2930_)
);

INV_X1 _7390_ (
  .A(_4557_),
  .ZN(_2931_)
);

XNOR2_X1 _7391_ (
  .A(_2930_),
  .B(_2931_),
  .ZN(_2932_)
);

AOI21_X1 _7392_ (
  .A(_2924_),
  .B1(_2932_),
  .B2(_1587_),
  .ZN(_0477_)
);

INV_X1 _7393_ (
  .A(_2920_),
  .ZN(_2933_)
);

NAND2_X1 _7394_ (
  .A1(_2922_),
  .A2(_4557_),
  .ZN(_2934_)
);

INV_X1 _7395_ (
  .A(_2934_),
  .ZN(_2935_)
);

NAND2_X1 _7396_ (
  .A1(_2933_),
  .A2(_2935_),
  .ZN(_2936_)
);

OR2_X2 _7397_ (
  .A1(_2906_),
  .A2(_2936_),
  .ZN(_2937_)
);

NAND2_X1 _7398_ (
  .A1(_2918_),
  .A2(_2935_),
  .ZN(_2938_)
);

INV_X1 _7399_ (
  .A(_4556_),
  .ZN(_2939_)
);

OAI21_X1 _7400_ (
  .A(_2939_),
  .B1(_2931_),
  .B2(_2925_),
  .ZN(_2940_)
);

INV_X1 _7401_ (
  .A(_2940_),
  .ZN(_2941_)
);

NAND2_X1 _7402_ (
  .A1(_2938_),
  .A2(_2941_),
  .ZN(_2942_)
);

INV_X1 _7403_ (
  .A(_2942_),
  .ZN(_2943_)
);

NAND2_X1 _7404_ (
  .A1(_2937_),
  .A2(_2943_),
  .ZN(_2944_)
);

NAND2_X1 _7405_ (
  .A1(_2944_),
  .A2(_4560_),
  .ZN(_2945_)
);

INV_X1 _7406_ (
  .A(_4560_),
  .ZN(_2946_)
);

NAND3_X1 _7407_ (
  .A1(_2937_),
  .A2(_2943_),
  .A3(_2946_),
  .ZN(_2947_)
);

NAND3_X1 _7408_ (
  .A1(_2945_),
  .A2(_2947_),
  .A3(_1572_),
  .ZN(_2948_)
);

INV_X1 _7409_ (
  .A(\s_pipe[5][19] ),
  .ZN(_2949_)
);

OAI21_X1 _7410_ (
  .A(_2948_),
  .B1(_2291_),
  .B2(_2949_),
  .ZN(_0478_)
);

NAND2_X1 _7411_ (
  .A1(_4557_),
  .A2(_4560_),
  .ZN(_2950_)
);

NOR2_X2 _7412_ (
  .A1(_2928_),
  .A2(_2950_),
  .ZN(_2951_)
);

NAND2_X1 _7413_ (
  .A1(_2912_),
  .A2(_2951_),
  .ZN(_2952_)
);

INV_X1 _7414_ (
  .A(_2950_),
  .ZN(_2953_)
);

NAND2_X1 _7415_ (
  .A1(_2927_),
  .A2(_2953_),
  .ZN(_2954_)
);

INV_X1 _7416_ (
  .A(_4559_),
  .ZN(_2955_)
);

OAI21_X1 _7417_ (
  .A(_2955_),
  .B1(_2946_),
  .B2(_2939_),
  .ZN(_2956_)
);

INV_X1 _7418_ (
  .A(_2956_),
  .ZN(_2957_)
);

NAND2_X1 _7419_ (
  .A1(_2954_),
  .A2(_2957_),
  .ZN(_2958_)
);

INV_X1 _7420_ (
  .A(_2958_),
  .ZN(_2959_)
);

NAND2_X1 _7421_ (
  .A1(_2952_),
  .A2(_2959_),
  .ZN(_2960_)
);

NAND2_X1 _7422_ (
  .A1(_2960_),
  .A2(_4563_),
  .ZN(_2961_)
);

INV_X1 _7423_ (
  .A(_4563_),
  .ZN(_2962_)
);

NAND3_X1 _7424_ (
  .A1(_2952_),
  .A2(_2959_),
  .A3(_2962_),
  .ZN(_2963_)
);

NAND3_X1 _7425_ (
  .A1(_2961_),
  .A2(_2963_),
  .A3(_1406_),
  .ZN(_2964_)
);

INV_X1 _7426_ (
  .A(\s_pipe[5][20] ),
  .ZN(_2965_)
);

OAI21_X1 _7427_ (
  .A(_2964_),
  .B1(_1351_),
  .B2(_2965_),
  .ZN(_0479_)
);

NAND2_X1 _7428_ (
  .A1(_2903_),
  .A2(_2933_),
  .ZN(_2966_)
);

NAND2_X1 _7429_ (
  .A1(_2966_),
  .A2(_2919_),
  .ZN(_2967_)
);

NAND2_X1 _7430_ (
  .A1(_4560_),
  .A2(_4563_),
  .ZN(_2968_)
);

NOR2_X1 _7431_ (
  .A1(_2934_),
  .A2(_2968_),
  .ZN(_2969_)
);

NAND2_X1 _7432_ (
  .A1(_2967_),
  .A2(_2969_),
  .ZN(_2970_)
);

INV_X1 _7433_ (
  .A(_2968_),
  .ZN(_2971_)
);

NAND2_X1 _7434_ (
  .A1(_2940_),
  .A2(_2971_),
  .ZN(_2972_)
);

INV_X1 _7435_ (
  .A(_4562_),
  .ZN(_2973_)
);

OAI21_X1 _7436_ (
  .A(_2973_),
  .B1(_2962_),
  .B2(_2955_),
  .ZN(_2974_)
);

INV_X1 _7437_ (
  .A(_2974_),
  .ZN(_2975_)
);

NAND2_X1 _7438_ (
  .A1(_2972_),
  .A2(_2975_),
  .ZN(_2976_)
);

INV_X1 _7439_ (
  .A(_2976_),
  .ZN(_2977_)
);

NOR2_X1 _7440_ (
  .A1(_2904_),
  .A2(_2920_),
  .ZN(_2978_)
);

NAND3_X1 _7441_ (
  .A1(_2978_),
  .A2(_2969_),
  .A3(_4121_),
  .ZN(_2979_)
);

NAND3_X1 _7442_ (
  .A1(_2970_),
  .A2(_2977_),
  .A3(_2979_),
  .ZN(_2980_)
);

NAND2_X1 _7443_ (
  .A1(_2980_),
  .A2(_4566_),
  .ZN(_2981_)
);

INV_X1 _7444_ (
  .A(_4566_),
  .ZN(_2982_)
);

NAND4_X1 _7445_ (
  .A1(_2970_),
  .A2(_2979_),
  .A3(_2977_),
  .A4(_2982_),
  .ZN(_2983_)
);

NAND3_X1 _7446_ (
  .A1(_2981_),
  .A2(_2983_),
  .A3(_1669_),
  .ZN(_2984_)
);

NAND2_X1 _7447_ (
  .A1(_1341_),
  .A2(\s_pipe[5][21] ),
  .ZN(_2985_)
);

NAND2_X1 _7448_ (
  .A1(_2984_),
  .A2(_2985_),
  .ZN(_0480_)
);

OAI21_X1 _7449_ (
  .A(_2911_),
  .B1(_2907_),
  .B2(_2901_),
  .ZN(_2986_)
);

NAND2_X1 _7450_ (
  .A1(_2986_),
  .A2(_2929_),
  .ZN(_2987_)
);

INV_X1 _7451_ (
  .A(_2927_),
  .ZN(_2988_)
);

NAND2_X1 _7452_ (
  .A1(_2987_),
  .A2(_2988_),
  .ZN(_2989_)
);

NAND2_X2 _7453_ (
  .A1(_4563_),
  .A2(_4566_),
  .ZN(_2990_)
);

NOR2_X1 _7454_ (
  .A1(_2950_),
  .A2(_2990_),
  .ZN(_2991_)
);

NAND2_X1 _7455_ (
  .A1(_2989_),
  .A2(_2991_),
  .ZN(_2992_)
);

INV_X2 _7456_ (
  .A(_2990_),
  .ZN(_2993_)
);

NAND2_X1 _7457_ (
  .A1(_2956_),
  .A2(_2993_),
  .ZN(_2994_)
);

INV_X1 _7458_ (
  .A(_4565_),
  .ZN(_2995_)
);

OAI21_X1 _7459_ (
  .A(_2995_),
  .B1(_2982_),
  .B2(_2973_),
  .ZN(_2996_)
);

INV_X1 _7460_ (
  .A(_2996_),
  .ZN(_2997_)
);

NAND2_X1 _7461_ (
  .A1(_2994_),
  .A2(_2997_),
  .ZN(_2998_)
);

INV_X1 _7462_ (
  .A(_2998_),
  .ZN(_2999_)
);

NOR3_X1 _7463_ (
  .A1(_2928_),
  .A2(_2896_),
  .A3(_2907_),
  .ZN(_3000_)
);

NAND3_X1 _7464_ (
  .A1(_3000_),
  .A2(_2991_),
  .A3(_2894_),
  .ZN(_3001_)
);

NAND3_X1 _7465_ (
  .A1(_2992_),
  .A2(_2999_),
  .A3(_3001_),
  .ZN(_3002_)
);

NAND2_X1 _7466_ (
  .A1(_3002_),
  .A2(_4569_),
  .ZN(_3003_)
);

INV_X1 _7467_ (
  .A(_4569_),
  .ZN(_3004_)
);

NAND4_X1 _7468_ (
  .A1(_2992_),
  .A2(_3001_),
  .A3(_2999_),
  .A4(_3004_),
  .ZN(_3005_)
);

NAND3_X1 _7469_ (
  .A1(_3003_),
  .A2(_3005_),
  .A3(_2001_),
  .ZN(_3006_)
);

NAND2_X1 _7470_ (
  .A1(_1709_),
  .A2(\s_pipe[5][22] ),
  .ZN(_3007_)
);

NAND2_X1 _7471_ (
  .A1(_3006_),
  .A2(_3007_),
  .ZN(_0481_)
);

NAND2_X1 _7472_ (
  .A1(_4566_),
  .A2(_4569_),
  .ZN(_3008_)
);

OR2_X2 _7473_ (
  .A1(_3008_),
  .A2(_2968_),
  .ZN(_3009_)
);

INV_X1 _7474_ (
  .A(_3009_),
  .ZN(_3010_)
);

NAND2_X1 _7475_ (
  .A1(_2942_),
  .A2(_3010_),
  .ZN(_3011_)
);

INV_X1 _7476_ (
  .A(_4568_),
  .ZN(_3012_)
);

OAI21_X1 _7477_ (
  .A(_3012_),
  .B1(_3004_),
  .B2(_2995_),
  .ZN(_3013_)
);

INV_X1 _7478_ (
  .A(_3013_),
  .ZN(_3014_)
);

OAI21_X1 _7479_ (
  .A(_3014_),
  .B1(_2975_),
  .B2(_3008_),
  .ZN(_3015_)
);

INV_X1 _7480_ (
  .A(_3015_),
  .ZN(_3016_)
);

INV_X1 _7481_ (
  .A(_2906_),
  .ZN(_3017_)
);

NOR2_X2 _7482_ (
  .A1(_3009_),
  .A2(_2936_),
  .ZN(_3018_)
);

NAND2_X1 _7483_ (
  .A1(_3017_),
  .A2(_3018_),
  .ZN(_3019_)
);

INV_X1 _7484_ (
  .A(_4572_),
  .ZN(_3020_)
);

NAND4_X1 _7485_ (
  .A1(_3011_),
  .A2(_3016_),
  .A3(_3019_),
  .A4(_3020_),
  .ZN(_3021_)
);

NAND3_X1 _7486_ (
  .A1(_3011_),
  .A2(_3016_),
  .A3(_3019_),
  .ZN(_3022_)
);

NAND2_X1 _7487_ (
  .A1(_3022_),
  .A2(_4572_),
  .ZN(_3023_)
);

NAND3_X1 _7488_ (
  .A1(_3021_),
  .A2(_3023_),
  .A3(_1669_),
  .ZN(_3024_)
);

NAND2_X1 _7489_ (
  .A1(_1341_),
  .A2(\s_pipe[5][23] ),
  .ZN(_3025_)
);

NAND2_X1 _7490_ (
  .A1(_3024_),
  .A2(_3025_),
  .ZN(_0482_)
);

NAND2_X1 _7491_ (
  .A1(_4569_),
  .A2(_4572_),
  .ZN(_3026_)
);

INV_X1 _7492_ (
  .A(_3026_),
  .ZN(_3027_)
);

NAND2_X1 _7493_ (
  .A1(_2993_),
  .A2(_3027_),
  .ZN(_3028_)
);

INV_X1 _7494_ (
  .A(_3028_),
  .ZN(_3029_)
);

NAND2_X1 _7495_ (
  .A1(_2958_),
  .A2(_3029_),
  .ZN(_3030_)
);

AND2_X2 _7496_ (
  .A1(_3029_),
  .A2(_2951_),
  .ZN(_3031_)
);

NAND2_X1 _7497_ (
  .A1(_2912_),
  .A2(_3031_),
  .ZN(_3032_)
);

NAND2_X1 _7498_ (
  .A1(_2996_),
  .A2(_3027_),
  .ZN(_3033_)
);

INV_X1 _7499_ (
  .A(_4571_),
  .ZN(_3034_)
);

OAI21_X1 _7500_ (
  .A(_3034_),
  .B1(_3020_),
  .B2(_3012_),
  .ZN(_3035_)
);

INV_X1 _7501_ (
  .A(_3035_),
  .ZN(_3036_)
);

NAND2_X1 _7502_ (
  .A1(_3033_),
  .A2(_3036_),
  .ZN(_3037_)
);

INV_X1 _7503_ (
  .A(_3037_),
  .ZN(_3038_)
);

NAND3_X2 _7504_ (
  .A1(_3030_),
  .A2(_3032_),
  .A3(_3038_),
  .ZN(_3039_)
);

INV_X1 _7505_ (
  .A(_3039_),
  .ZN(_3040_)
);

NOR2_X2 _7506_ (
  .A1(_1323_),
  .A2(\d_pipe[4][23] ),
  .ZN(_3041_)
);

NAND2_X4 _7507_ (
  .A1(_1307_),
  .A2(_3041_),
  .ZN(_3042_)
);

NAND2_X4 _7508_ (
  .A1(_3042_),
  .A2(_0657_),
  .ZN(_3043_)
);

INV_X1 _7509_ (
  .A(\s_pipe[4][23] ),
  .ZN(_3044_)
);

NAND2_X1 _7510_ (
  .A1(_3043_),
  .A2(_3044_),
  .ZN(_3045_)
);

NAND3_X1 _7511_ (
  .A1(_3042_),
  .A2(_0657_),
  .A3(\s_pipe[4][23] ),
  .ZN(_3046_)
);

NAND2_X1 _7512_ (
  .A1(_3045_),
  .A2(_3046_),
  .ZN(_3047_)
);

NAND2_X2 _7513_ (
  .A1(_3040_),
  .A2(_3047_),
  .ZN(_3048_)
);

NAND2_X1 _7514_ (
  .A1(_3043_),
  .A2(\s_pipe[4][23] ),
  .ZN(_3049_)
);

NAND3_X1 _7515_ (
  .A1(_3042_),
  .A2(_0657_),
  .A3(_3044_),
  .ZN(_3050_)
);

NAND2_X1 _7516_ (
  .A1(_3049_),
  .A2(_3050_),
  .ZN(_3051_)
);

NAND2_X1 _7517_ (
  .A1(_3051_),
  .A2(_3039_),
  .ZN(_3052_)
);

NAND3_X2 _7518_ (
  .A1(_3048_),
  .A2(_3052_),
  .A3(_1669_),
  .ZN(_3053_)
);

NAND2_X1 _7519_ (
  .A1(_1728_),
  .A2(\s_pipe[5][24] ),
  .ZN(_3054_)
);

NAND2_X2 _7520_ (
  .A1(_3053_),
  .A2(_3054_),
  .ZN(_0483_)
);

MUX2_X1 _7521_ (
  .A(\s_pipe[6][6] ),
  .B(\s_pipe[5][5] ),
  .S(_1566_),
  .Z(_0484_)
);

MUX2_X1 _7522_ (
  .A(\s_pipe[6][7] ),
  .B(\s_pipe[5][6] ),
  .S(_1563_),
  .Z(_0485_)
);

MUX2_X1 _7523_ (
  .A(\s_pipe[6][8] ),
  .B(\s_pipe[5][7] ),
  .S(_1563_),
  .Z(_0486_)
);

MUX2_X1 _7524_ (
  .A(\s_pipe[6][9] ),
  .B(\s_pipe[5][8] ),
  .S(_1563_),
  .Z(_0487_)
);

MUX2_X1 _7525_ (
  .A(\s_pipe[6][10] ),
  .B(\s_pipe[5][9] ),
  .S(_1563_),
  .Z(_0488_)
);

MUX2_X1 _7526_ (
  .A(\s_pipe[6][11] ),
  .B(\s_pipe[5][10] ),
  .S(_1563_),
  .Z(_0489_)
);

MUX2_X1 _7527_ (
  .A(\s_pipe[6][12] ),
  .B(_0127_),
  .S(_2068_),
  .Z(_0490_)
);

NAND2_X1 _7528_ (
  .A1(_1881_),
  .A2(\s_pipe[6][13] ),
  .ZN(_3055_)
);

OAI21_X1 _7529_ (
  .A(_3055_),
  .B1(_4112_),
  .B2(_2054_),
  .ZN(_0491_)
);

INV_X1 _7530_ (
  .A(_4111_),
  .ZN(_3056_)
);

NAND2_X1 _7531_ (
  .A1(_3056_),
  .A2(_4509_),
  .ZN(_3057_)
);

INV_X1 _7532_ (
  .A(_4509_),
  .ZN(_3058_)
);

NAND2_X1 _7533_ (
  .A1(_3058_),
  .A2(_4111_),
  .ZN(_3059_)
);

NAND3_X1 _7534_ (
  .A1(_3057_),
  .A2(_3059_),
  .A3(_1348_),
  .ZN(_3060_)
);

INV_X1 _7535_ (
  .A(\s_pipe[6][14] ),
  .ZN(_3061_)
);

OAI21_X1 _7536_ (
  .A(_3060_),
  .B1(_1634_),
  .B2(_3061_),
  .ZN(_0492_)
);

NOR2_X1 _7537_ (
  .A1(_1364_),
  .A2(\s_pipe[6][15] ),
  .ZN(_3062_)
);

INV_X1 _7538_ (
  .A(_4508_),
  .ZN(_3063_)
);

INV_X1 _7539_ (
  .A(_4505_),
  .ZN(_3064_)
);

OAI21_X1 _7540_ (
  .A(_3063_),
  .B1(_3058_),
  .B2(_3064_),
  .ZN(_3065_)
);

NAND2_X1 _7541_ (
  .A1(_4509_),
  .A2(_4506_),
  .ZN(_3066_)
);

NOR2_X1 _7542_ (
  .A1(_3066_),
  .A2(_4110_),
  .ZN(_3067_)
);

NOR2_X2 _7543_ (
  .A1(_3065_),
  .A2(_3067_),
  .ZN(_3068_)
);

INV_X1 _7544_ (
  .A(_4512_),
  .ZN(_3069_)
);

XNOR2_X1 _7545_ (
  .A(_3068_),
  .B(_3069_),
  .ZN(_3070_)
);

AOI21_X1 _7546_ (
  .A(_3062_),
  .B1(_3070_),
  .B2(_1901_),
  .ZN(_0493_)
);

NOR2_X1 _7547_ (
  .A1(_2091_),
  .A2(\s_pipe[6][16] ),
  .ZN(_3071_)
);

NOR2_X1 _7548_ (
  .A1(_4508_),
  .A2(_4511_),
  .ZN(_3072_)
);

INV_X1 _7549_ (
  .A(_4511_),
  .ZN(_3073_)
);

AOI22_X2 _7550_ (
  .A1(_3072_),
  .A2(_3057_),
  .B1(_3073_),
  .B2(_3069_),
  .ZN(_3074_)
);

BUF_X4 _7551_ (
  .A(_4515_),
  .Z(_3075_)
);

XNOR2_X1 _7552_ (
  .A(_3074_),
  .B(_3075_),
  .ZN(_3076_)
);

AOI21_X1 _7553_ (
  .A(_3071_),
  .B1(_3076_),
  .B2(_2265_),
  .ZN(_0494_)
);

NOR2_X1 _7554_ (
  .A1(_1371_),
  .A2(\s_pipe[6][17] ),
  .ZN(_3077_)
);

INV_X1 _7555_ (
  .A(_4514_),
  .ZN(_3078_)
);

INV_X1 _7556_ (
  .A(_3075_),
  .ZN(_3079_)
);

OAI21_X1 _7557_ (
  .A(_3078_),
  .B1(_3079_),
  .B2(_3073_),
  .ZN(_3080_)
);

INV_X1 _7558_ (
  .A(_3080_),
  .ZN(_3081_)
);

NAND2_X2 _7559_ (
  .A1(_4512_),
  .A2(_3075_),
  .ZN(_3082_)
);

OAI21_X1 _7560_ (
  .A(_3081_),
  .B1(_3068_),
  .B2(_3082_),
  .ZN(_3083_)
);

BUF_X4 _7561_ (
  .A(_4518_),
  .Z(_3084_)
);

XNOR2_X1 _7562_ (
  .A(_3083_),
  .B(_3084_),
  .ZN(_3085_)
);

AOI21_X1 _7563_ (
  .A(_3077_),
  .B1(_3085_),
  .B2(_1901_),
  .ZN(_0495_)
);

NOR2_X1 _7564_ (
  .A1(_1371_),
  .A2(\s_pipe[6][18] ),
  .ZN(_3086_)
);

INV_X1 _7565_ (
  .A(_4517_),
  .ZN(_3087_)
);

INV_X1 _7566_ (
  .A(_3084_),
  .ZN(_3088_)
);

OAI21_X2 _7567_ (
  .A(_3087_),
  .B1(_3088_),
  .B2(_3078_),
  .ZN(_3089_)
);

NAND2_X1 _7568_ (
  .A1(_3075_),
  .A2(_3084_),
  .ZN(_3090_)
);

INV_X1 _7569_ (
  .A(_3090_),
  .ZN(_3091_)
);

AOI21_X1 _7570_ (
  .A(_3089_),
  .B1(_3074_),
  .B2(_3091_),
  .ZN(_3092_)
);

INV_X1 _7571_ (
  .A(_4521_),
  .ZN(_3093_)
);

XNOR2_X1 _7572_ (
  .A(_3092_),
  .B(_3093_),
  .ZN(_3094_)
);

AOI21_X1 _7573_ (
  .A(_3086_),
  .B1(_3094_),
  .B2(_1587_),
  .ZN(_0496_)
);

INV_X1 _7574_ (
  .A(_3082_),
  .ZN(_3095_)
);

NAND2_X1 _7575_ (
  .A1(_3084_),
  .A2(_4521_),
  .ZN(_3096_)
);

INV_X1 _7576_ (
  .A(_3096_),
  .ZN(_3097_)
);

NAND2_X1 _7577_ (
  .A1(_3095_),
  .A2(_3097_),
  .ZN(_3098_)
);

OR2_X2 _7578_ (
  .A1(_3068_),
  .A2(_3098_),
  .ZN(_3099_)
);

NAND2_X1 _7579_ (
  .A1(_3080_),
  .A2(_3097_),
  .ZN(_3100_)
);

INV_X1 _7580_ (
  .A(_4520_),
  .ZN(_3101_)
);

OAI21_X1 _7581_ (
  .A(_3101_),
  .B1(_3093_),
  .B2(_3087_),
  .ZN(_3102_)
);

INV_X1 _7582_ (
  .A(_3102_),
  .ZN(_3103_)
);

NAND2_X1 _7583_ (
  .A1(_3100_),
  .A2(_3103_),
  .ZN(_3104_)
);

INV_X1 _7584_ (
  .A(_3104_),
  .ZN(_3105_)
);

NAND2_X1 _7585_ (
  .A1(_3099_),
  .A2(_3105_),
  .ZN(_3106_)
);

NAND2_X1 _7586_ (
  .A1(_3106_),
  .A2(_4524_),
  .ZN(_3107_)
);

INV_X1 _7587_ (
  .A(_4524_),
  .ZN(_3108_)
);

NAND3_X1 _7588_ (
  .A1(_3099_),
  .A2(_3105_),
  .A3(_3108_),
  .ZN(_3109_)
);

NAND3_X1 _7589_ (
  .A1(_3107_),
  .A2(_3109_),
  .A3(_2238_),
  .ZN(_3110_)
);

INV_X1 _7590_ (
  .A(\s_pipe[6][19] ),
  .ZN(_3111_)
);

OAI21_X1 _7591_ (
  .A(_3110_),
  .B1(_1901_),
  .B2(_3111_),
  .ZN(_0497_)
);

NAND2_X2 _7592_ (
  .A1(_4521_),
  .A2(_4524_),
  .ZN(_3112_)
);

NOR2_X2 _7593_ (
  .A1(_3090_),
  .A2(_3112_),
  .ZN(_3113_)
);

NAND2_X1 _7594_ (
  .A1(_3074_),
  .A2(_3113_),
  .ZN(_3114_)
);

INV_X1 _7595_ (
  .A(_3112_),
  .ZN(_3115_)
);

NAND2_X1 _7596_ (
  .A1(_3089_),
  .A2(_3115_),
  .ZN(_3116_)
);

INV_X1 _7597_ (
  .A(_4523_),
  .ZN(_3117_)
);

OAI21_X1 _7598_ (
  .A(_3117_),
  .B1(_3108_),
  .B2(_3101_),
  .ZN(_3118_)
);

INV_X1 _7599_ (
  .A(_3118_),
  .ZN(_3119_)
);

NAND2_X1 _7600_ (
  .A1(_3116_),
  .A2(_3119_),
  .ZN(_3120_)
);

INV_X1 _7601_ (
  .A(_3120_),
  .ZN(_3121_)
);

NAND2_X1 _7602_ (
  .A1(_3114_),
  .A2(_3121_),
  .ZN(_3122_)
);

NAND2_X1 _7603_ (
  .A1(_3122_),
  .A2(_4527_),
  .ZN(_3123_)
);

INV_X1 _7604_ (
  .A(_4527_),
  .ZN(_3124_)
);

NAND3_X1 _7605_ (
  .A1(_3114_),
  .A2(_3121_),
  .A3(_3124_),
  .ZN(_3125_)
);

NAND3_X1 _7606_ (
  .A1(_3123_),
  .A2(_3125_),
  .A3(_2238_),
  .ZN(_3126_)
);

INV_X1 _7607_ (
  .A(\s_pipe[6][20] ),
  .ZN(_3127_)
);

OAI21_X1 _7608_ (
  .A(_3126_),
  .B1(_1548_),
  .B2(_3127_),
  .ZN(_0498_)
);

NAND2_X1 _7609_ (
  .A1(_3065_),
  .A2(_3095_),
  .ZN(_3128_)
);

NAND2_X1 _7610_ (
  .A1(_3128_),
  .A2(_3081_),
  .ZN(_3129_)
);

NAND2_X2 _7611_ (
  .A1(_4524_),
  .A2(_4527_),
  .ZN(_3130_)
);

NOR2_X1 _7612_ (
  .A1(_3096_),
  .A2(_3130_),
  .ZN(_3131_)
);

NAND2_X1 _7613_ (
  .A1(_3129_),
  .A2(_3131_),
  .ZN(_3132_)
);

INV_X1 _7614_ (
  .A(_3130_),
  .ZN(_3133_)
);

NAND2_X1 _7615_ (
  .A1(_3102_),
  .A2(_3133_),
  .ZN(_3134_)
);

INV_X1 _7616_ (
  .A(_4526_),
  .ZN(_3135_)
);

OAI21_X1 _7617_ (
  .A(_3135_),
  .B1(_3124_),
  .B2(_3117_),
  .ZN(_3136_)
);

INV_X1 _7618_ (
  .A(_3136_),
  .ZN(_3137_)
);

NAND2_X1 _7619_ (
  .A1(_3134_),
  .A2(_3137_),
  .ZN(_3138_)
);

INV_X1 _7620_ (
  .A(_3138_),
  .ZN(_3139_)
);

NOR2_X1 _7621_ (
  .A1(_3066_),
  .A2(_3082_),
  .ZN(_3140_)
);

NAND3_X1 _7622_ (
  .A1(_3140_),
  .A2(_3131_),
  .A3(_4114_),
  .ZN(_3141_)
);

NAND3_X1 _7623_ (
  .A1(_3132_),
  .A2(_3139_),
  .A3(_3141_),
  .ZN(_3142_)
);

NAND2_X1 _7624_ (
  .A1(_3142_),
  .A2(_4530_),
  .ZN(_3143_)
);

INV_X1 _7625_ (
  .A(_4530_),
  .ZN(_3144_)
);

NAND4_X1 _7626_ (
  .A1(_3132_),
  .A2(_3141_),
  .A3(_3139_),
  .A4(_3144_),
  .ZN(_3145_)
);

NAND3_X1 _7627_ (
  .A1(_3143_),
  .A2(_3145_),
  .A3(_1447_),
  .ZN(_3146_)
);

NAND2_X1 _7628_ (
  .A1(_1341_),
  .A2(\s_pipe[6][21] ),
  .ZN(_3147_)
);

NAND2_X1 _7629_ (
  .A1(_3146_),
  .A2(_3147_),
  .ZN(_0499_)
);

OAI21_X1 _7630_ (
  .A(_3073_),
  .B1(_3069_),
  .B2(_3063_),
  .ZN(_3148_)
);

NAND2_X1 _7631_ (
  .A1(_3148_),
  .A2(_3091_),
  .ZN(_3149_)
);

INV_X1 _7632_ (
  .A(_3089_),
  .ZN(_3150_)
);

NAND2_X1 _7633_ (
  .A1(_3149_),
  .A2(_3150_),
  .ZN(_3151_)
);

NAND2_X2 _7634_ (
  .A1(_4527_),
  .A2(_4530_),
  .ZN(_3152_)
);

NOR2_X1 _7635_ (
  .A1(_3112_),
  .A2(_3152_),
  .ZN(_3153_)
);

NAND2_X1 _7636_ (
  .A1(_3151_),
  .A2(_3153_),
  .ZN(_3154_)
);

INV_X2 _7637_ (
  .A(_3152_),
  .ZN(_3155_)
);

NAND2_X1 _7638_ (
  .A1(_3118_),
  .A2(_3155_),
  .ZN(_3156_)
);

INV_X1 _7639_ (
  .A(_4529_),
  .ZN(_3157_)
);

OAI21_X1 _7640_ (
  .A(_3157_),
  .B1(_3144_),
  .B2(_3135_),
  .ZN(_3158_)
);

INV_X1 _7641_ (
  .A(_3158_),
  .ZN(_3159_)
);

NAND2_X1 _7642_ (
  .A1(_3156_),
  .A2(_3159_),
  .ZN(_3160_)
);

INV_X1 _7643_ (
  .A(_3160_),
  .ZN(_3161_)
);

NOR3_X1 _7644_ (
  .A1(_3090_),
  .A2(_3058_),
  .A3(_3069_),
  .ZN(_3162_)
);

NAND3_X1 _7645_ (
  .A1(_3162_),
  .A2(_3153_),
  .A3(_3056_),
  .ZN(_3163_)
);

NAND3_X1 _7646_ (
  .A1(_3154_),
  .A2(_3161_),
  .A3(_3163_),
  .ZN(_3164_)
);

NAND2_X1 _7647_ (
  .A1(_3164_),
  .A2(_4533_),
  .ZN(_3165_)
);

INV_X1 _7648_ (
  .A(_4533_),
  .ZN(_3166_)
);

NAND4_X1 _7649_ (
  .A1(_3154_),
  .A2(_3163_),
  .A3(_3161_),
  .A4(_3166_),
  .ZN(_3167_)
);

NAND3_X1 _7650_ (
  .A1(_3165_),
  .A2(_3167_),
  .A3(_1447_),
  .ZN(_3168_)
);

NAND2_X1 _7651_ (
  .A1(_1341_),
  .A2(\s_pipe[6][22] ),
  .ZN(_3169_)
);

NAND2_X1 _7652_ (
  .A1(_3168_),
  .A2(_3169_),
  .ZN(_0500_)
);

NAND2_X1 _7653_ (
  .A1(_4530_),
  .A2(_4533_),
  .ZN(_3170_)
);

OR2_X2 _7654_ (
  .A1(_3170_),
  .A2(_3130_),
  .ZN(_3171_)
);

INV_X1 _7655_ (
  .A(_3171_),
  .ZN(_3172_)
);

NAND2_X1 _7656_ (
  .A1(_3104_),
  .A2(_3172_),
  .ZN(_3173_)
);

INV_X1 _7657_ (
  .A(_4532_),
  .ZN(_3174_)
);

OAI21_X1 _7658_ (
  .A(_3174_),
  .B1(_3166_),
  .B2(_3157_),
  .ZN(_3175_)
);

INV_X1 _7659_ (
  .A(_3175_),
  .ZN(_3176_)
);

OAI21_X1 _7660_ (
  .A(_3176_),
  .B1(_3137_),
  .B2(_3170_),
  .ZN(_3177_)
);

INV_X1 _7661_ (
  .A(_3177_),
  .ZN(_3178_)
);

INV_X1 _7662_ (
  .A(_3068_),
  .ZN(_3179_)
);

NOR2_X2 _7663_ (
  .A1(_3171_),
  .A2(_3098_),
  .ZN(_3180_)
);

NAND2_X1 _7664_ (
  .A1(_3179_),
  .A2(_3180_),
  .ZN(_3181_)
);

INV_X1 _7665_ (
  .A(_4536_),
  .ZN(_3182_)
);

NAND4_X1 _7666_ (
  .A1(_3173_),
  .A2(_3178_),
  .A3(_3181_),
  .A4(_3182_),
  .ZN(_3183_)
);

NAND3_X1 _7667_ (
  .A1(_3173_),
  .A2(_3178_),
  .A3(_3181_),
  .ZN(_3184_)
);

NAND2_X1 _7668_ (
  .A1(_3184_),
  .A2(_4536_),
  .ZN(_3185_)
);

NAND3_X1 _7669_ (
  .A1(_3183_),
  .A2(_3185_),
  .A3(_2001_),
  .ZN(_3186_)
);

NAND2_X1 _7670_ (
  .A1(_1341_),
  .A2(\s_pipe[6][23] ),
  .ZN(_3187_)
);

NAND2_X1 _7671_ (
  .A1(_3186_),
  .A2(_3187_),
  .ZN(_0501_)
);

NAND2_X1 _7672_ (
  .A1(_4533_),
  .A2(_4536_),
  .ZN(_3188_)
);

INV_X1 _7673_ (
  .A(_3188_),
  .ZN(_3189_)
);

NAND2_X2 _7674_ (
  .A1(_3155_),
  .A2(_3189_),
  .ZN(_3190_)
);

INV_X2 _7675_ (
  .A(_3190_),
  .ZN(_3191_)
);

NAND2_X1 _7676_ (
  .A1(_3120_),
  .A2(_3191_),
  .ZN(_3192_)
);

AND2_X2 _7677_ (
  .A1(_3191_),
  .A2(_3113_),
  .ZN(_3193_)
);

NAND2_X2 _7678_ (
  .A1(_3074_),
  .A2(_3193_),
  .ZN(_3194_)
);

NAND2_X1 _7679_ (
  .A1(_3158_),
  .A2(_3189_),
  .ZN(_3195_)
);

INV_X1 _7680_ (
  .A(_4535_),
  .ZN(_3196_)
);

OAI21_X1 _7681_ (
  .A(_3196_),
  .B1(_3182_),
  .B2(_3174_),
  .ZN(_3197_)
);

INV_X1 _7682_ (
  .A(_3197_),
  .ZN(_3198_)
);

NAND2_X1 _7683_ (
  .A1(_3195_),
  .A2(_3198_),
  .ZN(_3199_)
);

INV_X1 _7684_ (
  .A(_3199_),
  .ZN(_3200_)
);

NAND3_X2 _7685_ (
  .A1(_3192_),
  .A2(_3194_),
  .A3(_3200_),
  .ZN(_3201_)
);

INV_X1 _7686_ (
  .A(_3201_),
  .ZN(_3202_)
);

NOR2_X2 _7687_ (
  .A1(_1260_),
  .A2(\d_pipe[5][23] ),
  .ZN(_3203_)
);

NAND2_X4 _7688_ (
  .A1(_1244_),
  .A2(_3203_),
  .ZN(_3204_)
);

NAND2_X4 _7689_ (
  .A1(_3204_),
  .A2(_0654_),
  .ZN(_3205_)
);

INV_X1 _7690_ (
  .A(\s_pipe[5][23] ),
  .ZN(_3206_)
);

NAND2_X1 _7691_ (
  .A1(_3205_),
  .A2(_3206_),
  .ZN(_3207_)
);

NAND3_X1 _7692_ (
  .A1(_3204_),
  .A2(_0654_),
  .A3(\s_pipe[5][23] ),
  .ZN(_3208_)
);

NAND2_X1 _7693_ (
  .A1(_3207_),
  .A2(_3208_),
  .ZN(_3209_)
);

NAND2_X1 _7694_ (
  .A1(_3202_),
  .A2(_3209_),
  .ZN(_3210_)
);

NAND2_X1 _7695_ (
  .A1(_3205_),
  .A2(\s_pipe[5][23] ),
  .ZN(_3211_)
);

NAND3_X1 _7696_ (
  .A1(_3204_),
  .A2(_0654_),
  .A3(_3206_),
  .ZN(_3212_)
);

NAND2_X1 _7697_ (
  .A1(_3211_),
  .A2(_3212_),
  .ZN(_3213_)
);

NAND2_X1 _7698_ (
  .A1(_3213_),
  .A2(_3201_),
  .ZN(_3214_)
);

NAND3_X1 _7699_ (
  .A1(_3210_),
  .A2(_3214_),
  .A3(_2001_),
  .ZN(_3215_)
);

NAND2_X1 _7700_ (
  .A1(_1341_),
  .A2(\s_pipe[6][24] ),
  .ZN(_3216_)
);

NAND2_X1 _7701_ (
  .A1(_3215_),
  .A2(_3216_),
  .ZN(_0502_)
);

NAND2_X1 _7702_ (
  .A1(_2349_),
  .A2(\s_pipe[9][9] ),
  .ZN(_3217_)
);

OAI21_X1 _7703_ (
  .A(_3217_),
  .B1(_1548_),
  .B2(_2400_),
  .ZN(_0503_)
);

MUX2_X1 _7704_ (
  .A(\s_pipe[10][11] ),
  .B(\s_pipe[9][10] ),
  .S(_1565_),
  .Z(_0504_)
);

MUX2_X1 _7705_ (
  .A(\s_pipe[10][12] ),
  .B(_0140_),
  .S(_1564_),
  .Z(_0505_)
);

NAND2_X1 _7706_ (
  .A1(_1338_),
  .A2(\s_pipe[10][13] ),
  .ZN(_3218_)
);

OAI21_X1 _7707_ (
  .A(_3218_),
  .B1(_4084_),
  .B2(_1562_),
  .ZN(_0506_)
);

INV_X1 _7708_ (
  .A(_4083_),
  .ZN(_3219_)
);

NAND2_X1 _7709_ (
  .A1(_3219_),
  .A2(_4365_),
  .ZN(_3220_)
);

INV_X1 _7710_ (
  .A(_4365_),
  .ZN(_3221_)
);

NAND2_X1 _7711_ (
  .A1(_3221_),
  .A2(_4083_),
  .ZN(_3222_)
);

NAND3_X1 _7712_ (
  .A1(_3220_),
  .A2(_3222_),
  .A3(_2238_),
  .ZN(_3223_)
);

INV_X1 _7713_ (
  .A(\s_pipe[10][14] ),
  .ZN(_3224_)
);

OAI21_X1 _7714_ (
  .A(_3223_),
  .B1(_2291_),
  .B2(_3224_),
  .ZN(_0507_)
);

NOR2_X1 _7715_ (
  .A1(_1371_),
  .A2(\s_pipe[10][15] ),
  .ZN(_3225_)
);

INV_X1 _7716_ (
  .A(_4364_),
  .ZN(_3226_)
);

INV_X1 _7717_ (
  .A(_4361_),
  .ZN(_3227_)
);

OAI21_X2 _7718_ (
  .A(_3226_),
  .B1(_3221_),
  .B2(_3227_),
  .ZN(_3228_)
);

NAND2_X1 _7719_ (
  .A1(_4365_),
  .A2(_4362_),
  .ZN(_3229_)
);

NOR2_X1 _7720_ (
  .A1(_3229_),
  .A2(_4082_),
  .ZN(_3230_)
);

NOR2_X2 _7721_ (
  .A1(_3228_),
  .A2(_3230_),
  .ZN(_3231_)
);

INV_X1 _7722_ (
  .A(_4368_),
  .ZN(_3232_)
);

XNOR2_X1 _7723_ (
  .A(_3231_),
  .B(_3232_),
  .ZN(_3233_)
);

AOI21_X1 _7724_ (
  .A(_3225_),
  .B1(_3233_),
  .B2(_1587_),
  .ZN(_0508_)
);

NOR2_X1 _7725_ (
  .A1(_1353_),
  .A2(\s_pipe[10][16] ),
  .ZN(_3234_)
);

NOR2_X1 _7726_ (
  .A1(_4364_),
  .A2(_4367_),
  .ZN(_3235_)
);

INV_X1 _7727_ (
  .A(_4367_),
  .ZN(_3236_)
);

AOI22_X2 _7728_ (
  .A1(_3235_),
  .A2(_3220_),
  .B1(_3236_),
  .B2(_3232_),
  .ZN(_3237_)
);

BUF_X4 _7729_ (
  .A(_4371_),
  .Z(_3238_)
);

XNOR2_X1 _7730_ (
  .A(_3237_),
  .B(_3238_),
  .ZN(_3239_)
);

AOI21_X1 _7731_ (
  .A(_3234_),
  .B1(_3239_),
  .B2(_1587_),
  .ZN(_0509_)
);

NOR2_X1 _7732_ (
  .A1(_1353_),
  .A2(\s_pipe[10][17] ),
  .ZN(_3240_)
);

INV_X1 _7733_ (
  .A(_4370_),
  .ZN(_3241_)
);

INV_X1 _7734_ (
  .A(_3238_),
  .ZN(_3242_)
);

OAI21_X1 _7735_ (
  .A(_3241_),
  .B1(_3242_),
  .B2(_3236_),
  .ZN(_3243_)
);

INV_X1 _7736_ (
  .A(_3243_),
  .ZN(_3244_)
);

NAND2_X2 _7737_ (
  .A1(_4368_),
  .A2(_3238_),
  .ZN(_3245_)
);

OAI21_X1 _7738_ (
  .A(_3244_),
  .B1(_3231_),
  .B2(_3245_),
  .ZN(_3246_)
);

BUF_X4 _7739_ (
  .A(_4374_),
  .Z(_3247_)
);

XNOR2_X1 _7740_ (
  .A(_3246_),
  .B(_3247_),
  .ZN(_3248_)
);

AOI21_X1 _7741_ (
  .A(_3240_),
  .B1(_3248_),
  .B2(_1587_),
  .ZN(_0510_)
);

NOR2_X1 _7742_ (
  .A1(_1364_),
  .A2(\s_pipe[10][18] ),
  .ZN(_3249_)
);

INV_X1 _7743_ (
  .A(_4373_),
  .ZN(_3250_)
);

INV_X1 _7744_ (
  .A(_3247_),
  .ZN(_3251_)
);

OAI21_X2 _7745_ (
  .A(_3250_),
  .B1(_3251_),
  .B2(_3241_),
  .ZN(_3252_)
);

NAND2_X1 _7746_ (
  .A1(_3238_),
  .A2(_3247_),
  .ZN(_3253_)
);

INV_X1 _7747_ (
  .A(_3253_),
  .ZN(_3254_)
);

AOI21_X1 _7748_ (
  .A(_3252_),
  .B1(_3237_),
  .B2(_3254_),
  .ZN(_3255_)
);

INV_X1 _7749_ (
  .A(_4377_),
  .ZN(_3256_)
);

XNOR2_X1 _7750_ (
  .A(_3255_),
  .B(_3256_),
  .ZN(_3257_)
);

AOI21_X1 _7751_ (
  .A(_3249_),
  .B1(_3257_),
  .B2(_1381_),
  .ZN(_0511_)
);

INV_X1 _7752_ (
  .A(_3245_),
  .ZN(_3258_)
);

NAND2_X1 _7753_ (
  .A1(_3247_),
  .A2(_4377_),
  .ZN(_3259_)
);

INV_X1 _7754_ (
  .A(_3259_),
  .ZN(_3260_)
);

NAND2_X1 _7755_ (
  .A1(_3258_),
  .A2(_3260_),
  .ZN(_3261_)
);

OR2_X2 _7756_ (
  .A1(_3231_),
  .A2(_3261_),
  .ZN(_3262_)
);

NAND2_X1 _7757_ (
  .A1(_3243_),
  .A2(_3260_),
  .ZN(_3263_)
);

INV_X1 _7758_ (
  .A(_4376_),
  .ZN(_3264_)
);

OAI21_X1 _7759_ (
  .A(_3264_),
  .B1(_3256_),
  .B2(_3250_),
  .ZN(_3265_)
);

INV_X1 _7760_ (
  .A(_3265_),
  .ZN(_3266_)
);

NAND2_X1 _7761_ (
  .A1(_3263_),
  .A2(_3266_),
  .ZN(_3267_)
);

INV_X1 _7762_ (
  .A(_3267_),
  .ZN(_3268_)
);

NAND2_X1 _7763_ (
  .A1(_3262_),
  .A2(_3268_),
  .ZN(_3269_)
);

NAND2_X1 _7764_ (
  .A1(_3269_),
  .A2(_4380_),
  .ZN(_3270_)
);

INV_X1 _7765_ (
  .A(_4380_),
  .ZN(_3271_)
);

NAND3_X1 _7766_ (
  .A1(_3262_),
  .A2(_3268_),
  .A3(_3271_),
  .ZN(_3272_)
);

NAND3_X1 _7767_ (
  .A1(_3270_),
  .A2(_3272_),
  .A3(_2238_),
  .ZN(_3273_)
);

INV_X1 _7768_ (
  .A(\s_pipe[10][19] ),
  .ZN(_3274_)
);

OAI21_X1 _7769_ (
  .A(_3273_),
  .B1(_1634_),
  .B2(_3274_),
  .ZN(_0512_)
);

NAND2_X1 _7770_ (
  .A1(_4377_),
  .A2(_4380_),
  .ZN(_3275_)
);

NOR2_X2 _7771_ (
  .A1(_3253_),
  .A2(_3275_),
  .ZN(_3276_)
);

NAND2_X1 _7772_ (
  .A1(_3237_),
  .A2(_3276_),
  .ZN(_3277_)
);

INV_X1 _7773_ (
  .A(_3275_),
  .ZN(_3278_)
);

NAND2_X1 _7774_ (
  .A1(_3252_),
  .A2(_3278_),
  .ZN(_3279_)
);

INV_X1 _7775_ (
  .A(_4379_),
  .ZN(_3280_)
);

OAI21_X1 _7776_ (
  .A(_3280_),
  .B1(_3271_),
  .B2(_3264_),
  .ZN(_3281_)
);

INV_X1 _7777_ (
  .A(_3281_),
  .ZN(_3282_)
);

NAND2_X1 _7778_ (
  .A1(_3279_),
  .A2(_3282_),
  .ZN(_3283_)
);

INV_X1 _7779_ (
  .A(_3283_),
  .ZN(_3284_)
);

NAND2_X1 _7780_ (
  .A1(_3277_),
  .A2(_3284_),
  .ZN(_3285_)
);

NAND2_X1 _7781_ (
  .A1(_3285_),
  .A2(_4383_),
  .ZN(_3286_)
);

INV_X1 _7782_ (
  .A(_4383_),
  .ZN(_3287_)
);

NAND3_X1 _7783_ (
  .A1(_3277_),
  .A2(_3284_),
  .A3(_3287_),
  .ZN(_3288_)
);

NAND3_X1 _7784_ (
  .A1(_3286_),
  .A2(_3288_),
  .A3(_2238_),
  .ZN(_3289_)
);

INV_X1 _7785_ (
  .A(\s_pipe[10][20] ),
  .ZN(_3290_)
);

OAI21_X1 _7786_ (
  .A(_3289_),
  .B1(_1408_),
  .B2(_3290_),
  .ZN(_0513_)
);

NAND2_X1 _7787_ (
  .A1(_3228_),
  .A2(_3258_),
  .ZN(_3291_)
);

NAND2_X1 _7788_ (
  .A1(_3291_),
  .A2(_3244_),
  .ZN(_3292_)
);

NAND2_X1 _7789_ (
  .A1(_4380_),
  .A2(_4383_),
  .ZN(_3293_)
);

NOR2_X1 _7790_ (
  .A1(_3259_),
  .A2(_3293_),
  .ZN(_3294_)
);

NAND2_X1 _7791_ (
  .A1(_3292_),
  .A2(_3294_),
  .ZN(_3295_)
);

INV_X1 _7792_ (
  .A(_3293_),
  .ZN(_3296_)
);

NAND2_X1 _7793_ (
  .A1(_3265_),
  .A2(_3296_),
  .ZN(_3297_)
);

INV_X1 _7794_ (
  .A(_4382_),
  .ZN(_3298_)
);

OAI21_X1 _7795_ (
  .A(_3298_),
  .B1(_3287_),
  .B2(_3280_),
  .ZN(_3299_)
);

INV_X1 _7796_ (
  .A(_3299_),
  .ZN(_3300_)
);

NAND2_X1 _7797_ (
  .A1(_3297_),
  .A2(_3300_),
  .ZN(_3301_)
);

INV_X1 _7798_ (
  .A(_3301_),
  .ZN(_3302_)
);

NOR2_X1 _7799_ (
  .A1(_3229_),
  .A2(_3245_),
  .ZN(_3303_)
);

NAND3_X1 _7800_ (
  .A1(_3303_),
  .A2(_3294_),
  .A3(_4086_),
  .ZN(_3304_)
);

NAND3_X1 _7801_ (
  .A1(_3295_),
  .A2(_3302_),
  .A3(_3304_),
  .ZN(_3305_)
);

NAND2_X1 _7802_ (
  .A1(_3305_),
  .A2(_4386_),
  .ZN(_3306_)
);

INV_X1 _7803_ (
  .A(_4386_),
  .ZN(_3307_)
);

NAND4_X1 _7804_ (
  .A1(_3295_),
  .A2(_3304_),
  .A3(_3302_),
  .A4(_3307_),
  .ZN(_3308_)
);

NAND3_X1 _7805_ (
  .A1(_3306_),
  .A2(_3308_),
  .A3(_2349_),
  .ZN(_3309_)
);

NAND2_X1 _7806_ (
  .A1(_1859_),
  .A2(\s_pipe[10][21] ),
  .ZN(_3310_)
);

NAND2_X1 _7807_ (
  .A1(_3309_),
  .A2(_3310_),
  .ZN(_0514_)
);

OAI21_X1 _7808_ (
  .A(_3236_),
  .B1(_3232_),
  .B2(_3226_),
  .ZN(_3311_)
);

NAND2_X1 _7809_ (
  .A1(_3311_),
  .A2(_3254_),
  .ZN(_3312_)
);

INV_X1 _7810_ (
  .A(_3252_),
  .ZN(_3313_)
);

NAND2_X1 _7811_ (
  .A1(_3312_),
  .A2(_3313_),
  .ZN(_3314_)
);

NAND2_X1 _7812_ (
  .A1(_4383_),
  .A2(_4386_),
  .ZN(_3315_)
);

NOR2_X1 _7813_ (
  .A1(_3275_),
  .A2(_3315_),
  .ZN(_3316_)
);

NAND2_X1 _7814_ (
  .A1(_3314_),
  .A2(_3316_),
  .ZN(_3317_)
);

INV_X2 _7815_ (
  .A(_3315_),
  .ZN(_3318_)
);

NAND2_X1 _7816_ (
  .A1(_3281_),
  .A2(_3318_),
  .ZN(_3319_)
);

INV_X1 _7817_ (
  .A(_4385_),
  .ZN(_3320_)
);

OAI21_X1 _7818_ (
  .A(_3320_),
  .B1(_3307_),
  .B2(_3298_),
  .ZN(_3321_)
);

INV_X1 _7819_ (
  .A(_3321_),
  .ZN(_3322_)
);

NAND2_X1 _7820_ (
  .A1(_3319_),
  .A2(_3322_),
  .ZN(_3323_)
);

INV_X1 _7821_ (
  .A(_3323_),
  .ZN(_3324_)
);

NOR3_X1 _7822_ (
  .A1(_3253_),
  .A2(_3221_),
  .A3(_3232_),
  .ZN(_3325_)
);

NAND3_X1 _7823_ (
  .A1(_3325_),
  .A2(_3316_),
  .A3(_3219_),
  .ZN(_3326_)
);

NAND3_X1 _7824_ (
  .A1(_3317_),
  .A2(_3324_),
  .A3(_3326_),
  .ZN(_3327_)
);

NAND2_X1 _7825_ (
  .A1(_3327_),
  .A2(_4389_),
  .ZN(_3328_)
);

INV_X1 _7826_ (
  .A(_4389_),
  .ZN(_3329_)
);

NAND4_X1 _7827_ (
  .A1(_3317_),
  .A2(_3326_),
  .A3(_3324_),
  .A4(_3329_),
  .ZN(_3330_)
);

NAND3_X1 _7828_ (
  .A1(_3328_),
  .A2(_3330_),
  .A3(_2001_),
  .ZN(_3331_)
);

NAND2_X1 _7829_ (
  .A1(_1859_),
  .A2(\s_pipe[10][22] ),
  .ZN(_3332_)
);

NAND2_X1 _7830_ (
  .A1(_3331_),
  .A2(_3332_),
  .ZN(_0515_)
);

NAND2_X1 _7831_ (
  .A1(_4386_),
  .A2(_4389_),
  .ZN(_3333_)
);

OR2_X2 _7832_ (
  .A1(_3333_),
  .A2(_3293_),
  .ZN(_3334_)
);

INV_X1 _7833_ (
  .A(_3334_),
  .ZN(_3335_)
);

NAND2_X1 _7834_ (
  .A1(_3267_),
  .A2(_3335_),
  .ZN(_3336_)
);

INV_X1 _7835_ (
  .A(_4388_),
  .ZN(_3337_)
);

OAI21_X1 _7836_ (
  .A(_3337_),
  .B1(_3329_),
  .B2(_3320_),
  .ZN(_3338_)
);

INV_X1 _7837_ (
  .A(_3338_),
  .ZN(_3339_)
);

OAI21_X1 _7838_ (
  .A(_3339_),
  .B1(_3300_),
  .B2(_3333_),
  .ZN(_3340_)
);

INV_X1 _7839_ (
  .A(_3340_),
  .ZN(_3341_)
);

INV_X1 _7840_ (
  .A(_3231_),
  .ZN(_3342_)
);

NOR2_X2 _7841_ (
  .A1(_3334_),
  .A2(_3261_),
  .ZN(_3343_)
);

NAND2_X1 _7842_ (
  .A1(_3342_),
  .A2(_3343_),
  .ZN(_3344_)
);

INV_X1 _7843_ (
  .A(_4392_),
  .ZN(_3345_)
);

NAND4_X1 _7844_ (
  .A1(_3336_),
  .A2(_3341_),
  .A3(_3344_),
  .A4(_3345_),
  .ZN(_3346_)
);

NAND3_X1 _7845_ (
  .A1(_3336_),
  .A2(_3341_),
  .A3(_3344_),
  .ZN(_3347_)
);

NAND2_X1 _7846_ (
  .A1(_3347_),
  .A2(_4392_),
  .ZN(_3348_)
);

NAND3_X1 _7847_ (
  .A1(_3346_),
  .A2(_3348_),
  .A3(_2001_),
  .ZN(_3349_)
);

NAND2_X1 _7848_ (
  .A1(_1859_),
  .A2(\s_pipe[10][23] ),
  .ZN(_3350_)
);

NAND2_X1 _7849_ (
  .A1(_3349_),
  .A2(_3350_),
  .ZN(_0516_)
);

NAND2_X1 _7850_ (
  .A1(_4389_),
  .A2(_4392_),
  .ZN(_3351_)
);

INV_X1 _7851_ (
  .A(_3351_),
  .ZN(_3352_)
);

NAND2_X2 _7852_ (
  .A1(_3318_),
  .A2(_3352_),
  .ZN(_3353_)
);

INV_X2 _7853_ (
  .A(_3353_),
  .ZN(_3354_)
);

NAND2_X1 _7854_ (
  .A1(_3283_),
  .A2(_3354_),
  .ZN(_3355_)
);

AND2_X2 _7855_ (
  .A1(_3354_),
  .A2(_3276_),
  .ZN(_3356_)
);

NAND2_X1 _7856_ (
  .A1(_3237_),
  .A2(_3356_),
  .ZN(_3357_)
);

NAND2_X1 _7857_ (
  .A1(_3321_),
  .A2(_3352_),
  .ZN(_3358_)
);

INV_X1 _7858_ (
  .A(_4391_),
  .ZN(_3359_)
);

OAI21_X1 _7859_ (
  .A(_3359_),
  .B1(_3345_),
  .B2(_3337_),
  .ZN(_3360_)
);

INV_X1 _7860_ (
  .A(_3360_),
  .ZN(_3361_)
);

NAND2_X1 _7861_ (
  .A1(_3358_),
  .A2(_3361_),
  .ZN(_3362_)
);

INV_X1 _7862_ (
  .A(_3362_),
  .ZN(_3363_)
);

NAND3_X2 _7863_ (
  .A1(_3355_),
  .A2(_3357_),
  .A3(_3363_),
  .ZN(_3364_)
);

INV_X1 _7864_ (
  .A(_3364_),
  .ZN(_3365_)
);

NOR2_X2 _7865_ (
  .A1(_1016_),
  .A2(_3713_),
  .ZN(_3366_)
);

NAND2_X4 _7866_ (
  .A1(_1001_),
  .A2(_3366_),
  .ZN(_3367_)
);

NAND2_X2 _7867_ (
  .A1(_3367_),
  .A2(_0642_),
  .ZN(_3368_)
);

INV_X1 _7868_ (
  .A(_0133_),
  .ZN(_3369_)
);

NAND2_X1 _7869_ (
  .A1(_3368_),
  .A2(_3369_),
  .ZN(_3370_)
);

NAND3_X1 _7870_ (
  .A1(_3367_),
  .A2(_0642_),
  .A3(_0133_),
  .ZN(_3371_)
);

NAND2_X1 _7871_ (
  .A1(_3370_),
  .A2(_3371_),
  .ZN(_3372_)
);

NAND2_X1 _7872_ (
  .A1(_3365_),
  .A2(_3372_),
  .ZN(_3373_)
);

NAND2_X1 _7873_ (
  .A1(_3368_),
  .A2(_0133_),
  .ZN(_3374_)
);

NAND3_X1 _7874_ (
  .A1(_3367_),
  .A2(_0642_),
  .A3(_3369_),
  .ZN(_3375_)
);

NAND2_X1 _7875_ (
  .A1(_3374_),
  .A2(_3375_),
  .ZN(_3376_)
);

NAND2_X1 _7876_ (
  .A1(_3376_),
  .A2(_3364_),
  .ZN(_3377_)
);

NAND3_X1 _7877_ (
  .A1(_3373_),
  .A2(_3377_),
  .A3(_1447_),
  .ZN(_3378_)
);

NAND2_X1 _7878_ (
  .A1(_1728_),
  .A2(\s_pipe[10][24] ),
  .ZN(_3379_)
);

NAND2_X1 _7879_ (
  .A1(_3378_),
  .A2(_3379_),
  .ZN(_0517_)
);

MUX2_X1 _7880_ (
  .A(\q_pipe[2][0] ),
  .B(_0112_),
  .S(_1861_),
  .Z(_0518_)
);

MUX2_X1 _7881_ (
  .A(\q_pipe[2][1] ),
  .B(\q_pipe[1] ),
  .S(_1861_),
  .Z(_0519_)
);

MUX2_X1 _7882_ (
  .A(\q_pipe[3][0] ),
  .B(_0113_),
  .S(_1934_),
  .Z(_0520_)
);

MUX2_X1 _7883_ (
  .A(\q_pipe[3][1] ),
  .B(\q_pipe[2][0] ),
  .S(_1934_),
  .Z(_0521_)
);

MUX2_X1 _7884_ (
  .A(\q_pipe[3][2] ),
  .B(\q_pipe[2][1] ),
  .S(_1861_),
  .Z(_0522_)
);

MUX2_X1 _7885_ (
  .A(\q_pipe[4][0] ),
  .B(_0114_),
  .S(_1952_),
  .Z(_0523_)
);

MUX2_X1 _7886_ (
  .A(\q_pipe[4][1] ),
  .B(\q_pipe[3][0] ),
  .S(_1861_),
  .Z(_0524_)
);

MUX2_X1 _7887_ (
  .A(\q_pipe[4][2] ),
  .B(\q_pipe[3][1] ),
  .S(_1861_),
  .Z(_0525_)
);

MUX2_X1 _7888_ (
  .A(\q_pipe[4][3] ),
  .B(\q_pipe[3][2] ),
  .S(_1861_),
  .Z(_0526_)
);

MUX2_X1 _7889_ (
  .A(\q_pipe[5][0] ),
  .B(_0115_),
  .S(_1566_),
  .Z(_0527_)
);

MUX2_X1 _7890_ (
  .A(\q_pipe[5][1] ),
  .B(\q_pipe[4][0] ),
  .S(_1566_),
  .Z(_0528_)
);

MUX2_X1 _7891_ (
  .A(\q_pipe[5][2] ),
  .B(\q_pipe[4][1] ),
  .S(_1566_),
  .Z(_0529_)
);

MUX2_X1 _7892_ (
  .A(\q_pipe[5][3] ),
  .B(\q_pipe[4][2] ),
  .S(_1566_),
  .Z(_0530_)
);

MUX2_X1 _7893_ (
  .A(\q_pipe[5][4] ),
  .B(\q_pipe[4][3] ),
  .S(_1566_),
  .Z(_0531_)
);

MUX2_X1 _7894_ (
  .A(\q_pipe[6][0] ),
  .B(_0116_),
  .S(_1563_),
  .Z(_0532_)
);

MUX2_X1 _7895_ (
  .A(\q_pipe[6][1] ),
  .B(\q_pipe[5][0] ),
  .S(_1563_),
  .Z(_0533_)
);

MUX2_X1 _7896_ (
  .A(\q_pipe[6][2] ),
  .B(\q_pipe[5][1] ),
  .S(_1563_),
  .Z(_0534_)
);

MUX2_X1 _7897_ (
  .A(\q_pipe[6][3] ),
  .B(\q_pipe[5][2] ),
  .S(_2007_),
  .Z(_0535_)
);

MUX2_X1 _7898_ (
  .A(\q_pipe[6][4] ),
  .B(\q_pipe[5][3] ),
  .S(_2007_),
  .Z(_0536_)
);

MUX2_X1 _7899_ (
  .A(\q_pipe[6][5] ),
  .B(\q_pipe[5][4] ),
  .S(_2007_),
  .Z(_0537_)
);

MUX2_X1 _7900_ (
  .A(\q_pipe[7][0] ),
  .B(_0117_),
  .S(_1952_),
  .Z(_0538_)
);

MUX2_X1 _7901_ (
  .A(\q_pipe[7][1] ),
  .B(\q_pipe[6][0] ),
  .S(_1952_),
  .Z(_0539_)
);

MUX2_X1 _7902_ (
  .A(\q_pipe[7][2] ),
  .B(\q_pipe[6][1] ),
  .S(_1952_),
  .Z(_0540_)
);

MUX2_X1 _7903_ (
  .A(\q_pipe[7][3] ),
  .B(\q_pipe[6][2] ),
  .S(_1952_),
  .Z(_0541_)
);

MUX2_X1 _7904_ (
  .A(\q_pipe[7][4] ),
  .B(\q_pipe[6][3] ),
  .S(_1952_),
  .Z(_0542_)
);

MUX2_X1 _7905_ (
  .A(\q_pipe[7][5] ),
  .B(\q_pipe[6][4] ),
  .S(_2068_),
  .Z(_0543_)
);

MUX2_X1 _7906_ (
  .A(\q_pipe[7][6] ),
  .B(\q_pipe[6][5] ),
  .S(_2068_),
  .Z(_0544_)
);

MUX2_X1 _7907_ (
  .A(\q_pipe[8][0] ),
  .B(_0118_),
  .S(_2068_),
  .Z(_0545_)
);

MUX2_X1 _7908_ (
  .A(\q_pipe[8][1] ),
  .B(\q_pipe[7][0] ),
  .S(_2068_),
  .Z(_0546_)
);

MUX2_X1 _7909_ (
  .A(\q_pipe[8][2] ),
  .B(\q_pipe[7][1] ),
  .S(_2068_),
  .Z(_0547_)
);

MUX2_X1 _7910_ (
  .A(\q_pipe[8][3] ),
  .B(\q_pipe[7][2] ),
  .S(_2067_),
  .Z(_0548_)
);

MUX2_X1 _7911_ (
  .A(\q_pipe[8][4] ),
  .B(\q_pipe[7][3] ),
  .S(_2067_),
  .Z(_0549_)
);

MUX2_X1 _7912_ (
  .A(\q_pipe[8][5] ),
  .B(\q_pipe[7][4] ),
  .S(_2067_),
  .Z(_0550_)
);

MUX2_X1 _7913_ (
  .A(\q_pipe[8][6] ),
  .B(\q_pipe[7][5] ),
  .S(_2067_),
  .Z(_0551_)
);

MUX2_X1 _7914_ (
  .A(\q_pipe[8][7] ),
  .B(\q_pipe[7][6] ),
  .S(_2067_),
  .Z(_0552_)
);

MUX2_X1 _7915_ (
  .A(\q_pipe[9] ),
  .B(_0119_),
  .S(_2067_),
  .Z(_0553_)
);

MUX2_X1 _7916_ (
  .A(_0618_),
  .B(\q_pipe[8][0] ),
  .S(_1898_),
  .Z(_0554_)
);

MUX2_X1 _7917_ (
  .A(_0619_),
  .B(\q_pipe[8][1] ),
  .S(_1898_),
  .Z(_0555_)
);

MUX2_X1 _7918_ (
  .A(_0620_),
  .B(\q_pipe[8][2] ),
  .S(_1897_),
  .Z(_0556_)
);

MUX2_X1 _7919_ (
  .A(_0621_),
  .B(\q_pipe[8][3] ),
  .S(_1897_),
  .Z(_0557_)
);

MUX2_X1 _7920_ (
  .A(_0622_),
  .B(\q_pipe[8][4] ),
  .S(_2066_),
  .Z(_0558_)
);

MUX2_X1 _7921_ (
  .A(_0623_),
  .B(\q_pipe[8][5] ),
  .S(_2066_),
  .Z(_0559_)
);

MUX2_X1 _7922_ (
  .A(_0624_),
  .B(\q_pipe[8][6] ),
  .S(_2066_),
  .Z(_0560_)
);

MUX2_X1 _7923_ (
  .A(_0625_),
  .B(\q_pipe[8][7] ),
  .S(_2066_),
  .Z(_0561_)
);

MUX2_X1 _7924_ (
  .A(\q_pipe[10][0] ),
  .B(_0120_),
  .S(_2066_),
  .Z(_0562_)
);

MUX2_X1 _7925_ (
  .A(\q_pipe[10][1] ),
  .B(\q_pipe[9] ),
  .S(_2066_),
  .Z(_0563_)
);

MUX2_X1 _7926_ (
  .A(\q_pipe[10][2] ),
  .B(_0618_),
  .S(_1565_),
  .Z(_0564_)
);

MUX2_X1 _7927_ (
  .A(\q_pipe[10][3] ),
  .B(_0619_),
  .S(_1565_),
  .Z(_0565_)
);

MUX2_X1 _7928_ (
  .A(\q_pipe[10][4] ),
  .B(_0620_),
  .S(_1564_),
  .Z(_0566_)
);

MUX2_X1 _7929_ (
  .A(\q_pipe[10][5] ),
  .B(_0621_),
  .S(_1564_),
  .Z(_0567_)
);

MUX2_X1 _7930_ (
  .A(\q_pipe[10][6] ),
  .B(_0622_),
  .S(_2007_),
  .Z(_0568_)
);

MUX2_X1 _7931_ (
  .A(\q_pipe[10][7] ),
  .B(_0623_),
  .S(_2007_),
  .Z(_0569_)
);

MUX2_X1 _7932_ (
  .A(\q_pipe[10][8] ),
  .B(_0624_),
  .S(_1933_),
  .Z(_0570_)
);

MUX2_X1 _7933_ (
  .A(\q_pipe[10][9] ),
  .B(_0625_),
  .S(_1933_),
  .Z(_0571_)
);

NAND2_X1 _7934_ (
  .A1(_1546_),
  .A2(_0121_),
  .ZN(_3380_)
);

OAI21_X1 _7935_ (
  .A(_3380_),
  .B1(_2291_),
  .B2(_1863_),
  .ZN(_0572_)
);

NAND2_X1 _7936_ (
  .A1(_1899_),
  .A2(\q_pipe[10][0] ),
  .ZN(_3381_)
);

OAI21_X1 _7937_ (
  .A(_3381_),
  .B1(_2291_),
  .B2(_1866_),
  .ZN(_0573_)
);

NAND2_X1 _7938_ (
  .A1(_1899_),
  .A2(\q_pipe[10][1] ),
  .ZN(_3382_)
);

OAI21_X1 _7939_ (
  .A(_3382_),
  .B1(_2291_),
  .B2(_1868_),
  .ZN(_0574_)
);

NAND2_X1 _7940_ (
  .A1(_1899_),
  .A2(\q_pipe[10][2] ),
  .ZN(_3383_)
);

OAI21_X1 _7941_ (
  .A(_3383_),
  .B1(_1548_),
  .B2(_1870_),
  .ZN(_0575_)
);

NAND2_X1 _7942_ (
  .A1(_1899_),
  .A2(\q_pipe[10][3] ),
  .ZN(_3384_)
);

OAI21_X1 _7943_ (
  .A(_3384_),
  .B1(_1548_),
  .B2(_1872_),
  .ZN(_0576_)
);

NAND2_X1 _7944_ (
  .A1(_1899_),
  .A2(\q_pipe[10][4] ),
  .ZN(_3385_)
);

OAI21_X1 _7945_ (
  .A(_3385_),
  .B1(_1901_),
  .B2(_1874_),
  .ZN(_0577_)
);

NAND2_X1 _7946_ (
  .A1(_1899_),
  .A2(\q_pipe[10][5] ),
  .ZN(_3386_)
);

OAI21_X1 _7947_ (
  .A(_3386_),
  .B1(_1548_),
  .B2(_1876_),
  .ZN(_0578_)
);

NAND2_X1 _7948_ (
  .A1(_1899_),
  .A2(\q_pipe[10][6] ),
  .ZN(_3387_)
);

OAI21_X1 _7949_ (
  .A(_3387_),
  .B1(_1408_),
  .B2(_1878_),
  .ZN(_0579_)
);

NAND2_X1 _7950_ (
  .A1(_1899_),
  .A2(\q_pipe[10][7] ),
  .ZN(_3388_)
);

OAI21_X1 _7951_ (
  .A(_3388_),
  .B1(_1634_),
  .B2(_1880_),
  .ZN(_0580_)
);

NAND2_X1 _7952_ (
  .A1(_1546_),
  .A2(\q_pipe[10][8] ),
  .ZN(_3389_)
);

OAI21_X1 _7953_ (
  .A(_3389_),
  .B1(_1634_),
  .B2(_1883_),
  .ZN(_0581_)
);

NAND2_X1 _7954_ (
  .A1(_2349_),
  .A2(\q_pipe[10][9] ),
  .ZN(_3390_)
);

OAI21_X1 _7955_ (
  .A(_3390_),
  .B1(_1634_),
  .B2(_1885_),
  .ZN(_0582_)
);

MUX2_X1 _7956_ (
  .A(\s_pipe[7][7] ),
  .B(\s_pipe[6][6] ),
  .S(_1897_),
  .Z(_0583_)
);

MUX2_X1 _7957_ (
  .A(\s_pipe[7][8] ),
  .B(\s_pipe[6][7] ),
  .S(_1897_),
  .Z(_0584_)
);

MUX2_X1 _7958_ (
  .A(\s_pipe[7][9] ),
  .B(\s_pipe[6][8] ),
  .S(_1897_),
  .Z(_0585_)
);

MUX2_X1 _7959_ (
  .A(\s_pipe[7][10] ),
  .B(\s_pipe[6][9] ),
  .S(_1897_),
  .Z(_0586_)
);

MUX2_X1 _7960_ (
  .A(\s_pipe[7][11] ),
  .B(\s_pipe[6][10] ),
  .S(_1934_),
  .Z(_0587_)
);

MUX2_X1 _7961_ (
  .A(\s_pipe[7][12] ),
  .B(_0128_),
  .S(_1934_),
  .Z(_0588_)
);

NAND2_X1 _7962_ (
  .A1(_1522_),
  .A2(\s_pipe[7][13] ),
  .ZN(_3391_)
);

OAI21_X1 _7963_ (
  .A(_3391_),
  .B1(_4105_),
  .B2(_1562_),
  .ZN(_0589_)
);

INV_X1 _7964_ (
  .A(_4104_),
  .ZN(_3392_)
);

NAND2_X1 _7965_ (
  .A1(_3392_),
  .A2(_4473_),
  .ZN(_3393_)
);

INV_X2 _7966_ (
  .A(_4473_),
  .ZN(_3394_)
);

NAND2_X1 _7967_ (
  .A1(_3394_),
  .A2(_4104_),
  .ZN(_3395_)
);

NAND3_X1 _7968_ (
  .A1(_3393_),
  .A2(_3395_),
  .A3(_1348_),
  .ZN(_3396_)
);

INV_X1 _7969_ (
  .A(\s_pipe[7][14] ),
  .ZN(_3397_)
);

OAI21_X1 _7970_ (
  .A(_3396_),
  .B1(_1901_),
  .B2(_3397_),
  .ZN(_0590_)
);

NOR2_X1 _7971_ (
  .A1(_1364_),
  .A2(\s_pipe[7][15] ),
  .ZN(_3398_)
);

INV_X1 _7972_ (
  .A(_4472_),
  .ZN(_3399_)
);

INV_X1 _7973_ (
  .A(_4469_),
  .ZN(_3400_)
);

OAI21_X1 _7974_ (
  .A(_3399_),
  .B1(_3394_),
  .B2(_3400_),
  .ZN(_3401_)
);

NAND2_X1 _7975_ (
  .A1(_4473_),
  .A2(_4470_),
  .ZN(_3402_)
);

NOR2_X1 _7976_ (
  .A1(_3402_),
  .A2(_4103_),
  .ZN(_3403_)
);

NOR2_X2 _7977_ (
  .A1(_3401_),
  .A2(_3403_),
  .ZN(_3404_)
);

INV_X1 _7978_ (
  .A(_4476_),
  .ZN(_3405_)
);

XNOR2_X1 _7979_ (
  .A(_3404_),
  .B(_3405_),
  .ZN(_3406_)
);

AOI21_X1 _7980_ (
  .A(_3398_),
  .B1(_3406_),
  .B2(_1552_),
  .ZN(_0591_)
);

NOR2_X1 _7981_ (
  .A1(_1371_),
  .A2(\s_pipe[7][16] ),
  .ZN(_3407_)
);

INV_X1 _7982_ (
  .A(_4475_),
  .ZN(_3408_)
);

OAI21_X2 _7983_ (
  .A(_3408_),
  .B1(_3405_),
  .B2(_3399_),
  .ZN(_3409_)
);

INV_X2 _7984_ (
  .A(_3409_),
  .ZN(_3410_)
);

NAND3_X1 _7985_ (
  .A1(_3392_),
  .A2(_4473_),
  .A3(_4476_),
  .ZN(_3411_)
);

NAND2_X2 _7986_ (
  .A1(_3410_),
  .A2(_3411_),
  .ZN(_3412_)
);

BUF_X2 _7987_ (
  .A(_4479_),
  .Z(_3413_)
);

XNOR2_X1 _7988_ (
  .A(_3412_),
  .B(_3413_),
  .ZN(_3414_)
);

AOI21_X1 _7989_ (
  .A(_3407_),
  .B1(_3414_),
  .B2(_1381_),
  .ZN(_0592_)
);

NOR2_X1 _7990_ (
  .A1(_1364_),
  .A2(\s_pipe[7][17] ),
  .ZN(_3415_)
);

INV_X1 _7991_ (
  .A(_4478_),
  .ZN(_3416_)
);

INV_X1 _7992_ (
  .A(_3413_),
  .ZN(_3417_)
);

OAI21_X1 _7993_ (
  .A(_3416_),
  .B1(_3417_),
  .B2(_3408_),
  .ZN(_3418_)
);

INV_X1 _7994_ (
  .A(_3418_),
  .ZN(_3419_)
);

NAND2_X2 _7995_ (
  .A1(_4476_),
  .A2(_3413_),
  .ZN(_3420_)
);

OAI21_X2 _7996_ (
  .A(_3419_),
  .B1(_3404_),
  .B2(_3420_),
  .ZN(_3421_)
);

BUF_X4 _7997_ (
  .A(_4482_),
  .Z(_3422_)
);

XNOR2_X1 _7998_ (
  .A(_3421_),
  .B(_3422_),
  .ZN(_3423_)
);

AOI21_X1 _7999_ (
  .A(_3415_),
  .B1(_3423_),
  .B2(_1381_),
  .ZN(_0593_)
);

NOR2_X1 _8000_ (
  .A1(_1353_),
  .A2(\s_pipe[7][18] ),
  .ZN(_3424_)
);

NAND2_X2 _8001_ (
  .A1(_3422_),
  .A2(_4478_),
  .ZN(_3425_)
);

INV_X1 _8002_ (
  .A(_4481_),
  .ZN(_3426_)
);

NAND2_X2 _8003_ (
  .A1(_3425_),
  .A2(_3426_),
  .ZN(_3427_)
);

NAND2_X2 _8004_ (
  .A1(_3413_),
  .A2(_3422_),
  .ZN(_3428_)
);

INV_X1 _8005_ (
  .A(_3428_),
  .ZN(_3429_)
);

AOI21_X2 _8006_ (
  .A(_3427_),
  .B1(_3412_),
  .B2(_3429_),
  .ZN(_3430_)
);

INV_X1 _8007_ (
  .A(_4485_),
  .ZN(_3431_)
);

XNOR2_X1 _8008_ (
  .A(_3430_),
  .B(_3431_),
  .ZN(_3432_)
);

AOI21_X1 _8009_ (
  .A(_3424_),
  .B1(_3432_),
  .B2(_1587_),
  .ZN(_0594_)
);

INV_X2 _8010_ (
  .A(_3420_),
  .ZN(_3433_)
);

NAND2_X1 _8011_ (
  .A1(_3422_),
  .A2(_4485_),
  .ZN(_3434_)
);

INV_X1 _8012_ (
  .A(_3434_),
  .ZN(_3435_)
);

NAND2_X1 _8013_ (
  .A1(_3433_),
  .A2(_3435_),
  .ZN(_3436_)
);

OR2_X2 _8014_ (
  .A1(_3404_),
  .A2(_3436_),
  .ZN(_3437_)
);

NAND2_X1 _8015_ (
  .A1(_3418_),
  .A2(_3435_),
  .ZN(_3438_)
);

INV_X1 _8016_ (
  .A(_4484_),
  .ZN(_3439_)
);

OAI21_X1 _8017_ (
  .A(_3439_),
  .B1(_3431_),
  .B2(_3426_),
  .ZN(_3440_)
);

INV_X1 _8018_ (
  .A(_3440_),
  .ZN(_3441_)
);

NAND2_X1 _8019_ (
  .A1(_3438_),
  .A2(_3441_),
  .ZN(_3442_)
);

INV_X1 _8020_ (
  .A(_3442_),
  .ZN(_3443_)
);

NAND2_X1 _8021_ (
  .A1(_3437_),
  .A2(_3443_),
  .ZN(_3444_)
);

NAND2_X1 _8022_ (
  .A1(_3444_),
  .A2(_4488_),
  .ZN(_3445_)
);

INV_X1 _8023_ (
  .A(_4488_),
  .ZN(_3446_)
);

NAND3_X1 _8024_ (
  .A1(_3437_),
  .A2(_3443_),
  .A3(_3446_),
  .ZN(_3447_)
);

NAND3_X1 _8025_ (
  .A1(_3445_),
  .A2(_3447_),
  .A3(_1572_),
  .ZN(_3448_)
);

INV_X1 _8026_ (
  .A(\s_pipe[7][19] ),
  .ZN(_3449_)
);

OAI21_X1 _8027_ (
  .A(_3448_),
  .B1(_1351_),
  .B2(_3449_),
  .ZN(_0595_)
);

NAND2_X1 _8028_ (
  .A1(_4485_),
  .A2(_4488_),
  .ZN(_3450_)
);

NOR2_X2 _8029_ (
  .A1(_3428_),
  .A2(_3450_),
  .ZN(_3451_)
);

NAND2_X1 _8030_ (
  .A1(_3412_),
  .A2(_3451_),
  .ZN(_3452_)
);

INV_X1 _8031_ (
  .A(_4487_),
  .ZN(_3453_)
);

OAI21_X1 _8032_ (
  .A(_3453_),
  .B1(_3446_),
  .B2(_3439_),
  .ZN(_3454_)
);

INV_X1 _8033_ (
  .A(_3454_),
  .ZN(_3455_)
);

INV_X1 _8034_ (
  .A(_3450_),
  .ZN(_3456_)
);

NAND2_X1 _8035_ (
  .A1(_3427_),
  .A2(_3456_),
  .ZN(_3457_)
);

NAND2_X1 _8036_ (
  .A1(_3455_),
  .A2(_3457_),
  .ZN(_3458_)
);

INV_X1 _8037_ (
  .A(_3458_),
  .ZN(_3459_)
);

NAND2_X1 _8038_ (
  .A1(_3452_),
  .A2(_3459_),
  .ZN(_3460_)
);

NAND2_X1 _8039_ (
  .A1(_3460_),
  .A2(_4491_),
  .ZN(_3461_)
);

INV_X1 _8040_ (
  .A(_4491_),
  .ZN(_3462_)
);

NAND3_X1 _8041_ (
  .A1(_3452_),
  .A2(_3462_),
  .A3(_3459_),
  .ZN(_3463_)
);

NAND3_X1 _8042_ (
  .A1(_3461_),
  .A2(_3463_),
  .A3(_1572_),
  .ZN(_3464_)
);

INV_X1 _8043_ (
  .A(\s_pipe[7][20] ),
  .ZN(_3465_)
);

OAI21_X1 _8044_ (
  .A(_3464_),
  .B1(_1351_),
  .B2(_3465_),
  .ZN(_0596_)
);

NAND2_X1 _8045_ (
  .A1(_3401_),
  .A2(_3433_),
  .ZN(_3466_)
);

NAND2_X1 _8046_ (
  .A1(_3466_),
  .A2(_3419_),
  .ZN(_3467_)
);

NAND2_X1 _8047_ (
  .A1(_4488_),
  .A2(_4491_),
  .ZN(_3468_)
);

NOR2_X1 _8048_ (
  .A1(_3434_),
  .A2(_3468_),
  .ZN(_3469_)
);

NAND2_X1 _8049_ (
  .A1(_3467_),
  .A2(_3469_),
  .ZN(_3470_)
);

INV_X1 _8050_ (
  .A(_3468_),
  .ZN(_3471_)
);

NAND2_X1 _8051_ (
  .A1(_3440_),
  .A2(_3471_),
  .ZN(_3472_)
);

INV_X1 _8052_ (
  .A(_4490_),
  .ZN(_3473_)
);

OAI21_X1 _8053_ (
  .A(_3473_),
  .B1(_3462_),
  .B2(_3453_),
  .ZN(_3474_)
);

INV_X1 _8054_ (
  .A(_3474_),
  .ZN(_3475_)
);

NAND2_X1 _8055_ (
  .A1(_3472_),
  .A2(_3475_),
  .ZN(_3476_)
);

INV_X1 _8056_ (
  .A(_3476_),
  .ZN(_3477_)
);

NOR2_X1 _8057_ (
  .A1(_3402_),
  .A2(_3420_),
  .ZN(_3478_)
);

NAND3_X1 _8058_ (
  .A1(_3478_),
  .A2(_3469_),
  .A3(_4107_),
  .ZN(_3479_)
);

NAND3_X1 _8059_ (
  .A1(_3470_),
  .A2(_3477_),
  .A3(_3479_),
  .ZN(_3480_)
);

NAND2_X1 _8060_ (
  .A1(_3480_),
  .A2(_4494_),
  .ZN(_3481_)
);

INV_X1 _8061_ (
  .A(_4494_),
  .ZN(_3482_)
);

NAND4_X1 _8062_ (
  .A1(_3470_),
  .A2(_3479_),
  .A3(_3477_),
  .A4(_3482_),
  .ZN(_3483_)
);

NAND3_X1 _8063_ (
  .A1(_3481_),
  .A2(_3483_),
  .A3(_1669_),
  .ZN(_3484_)
);

NAND2_X1 _8064_ (
  .A1(_1728_),
  .A2(\s_pipe[7][21] ),
  .ZN(_3485_)
);

NAND2_X1 _8065_ (
  .A1(_3484_),
  .A2(_3485_),
  .ZN(_0597_)
);

NAND2_X1 _8066_ (
  .A1(_3409_),
  .A2(_3429_),
  .ZN(_3486_)
);

INV_X1 _8067_ (
  .A(_3427_),
  .ZN(_3487_)
);

NAND2_X1 _8068_ (
  .A1(_3486_),
  .A2(_3487_),
  .ZN(_3488_)
);

NAND2_X1 _8069_ (
  .A1(_4491_),
  .A2(_4494_),
  .ZN(_3489_)
);

NOR2_X1 _8070_ (
  .A1(_3450_),
  .A2(_3489_),
  .ZN(_3490_)
);

NAND2_X1 _8071_ (
  .A1(_3488_),
  .A2(_3490_),
  .ZN(_3491_)
);

INV_X1 _8072_ (
  .A(_3489_),
  .ZN(_3492_)
);

NAND2_X1 _8073_ (
  .A1(_3454_),
  .A2(_3492_),
  .ZN(_3493_)
);

INV_X1 _8074_ (
  .A(_4493_),
  .ZN(_3494_)
);

OAI21_X1 _8075_ (
  .A(_3494_),
  .B1(_3482_),
  .B2(_3473_),
  .ZN(_3495_)
);

INV_X1 _8076_ (
  .A(_3495_),
  .ZN(_3496_)
);

NAND2_X1 _8077_ (
  .A1(_3493_),
  .A2(_3496_),
  .ZN(_3497_)
);

INV_X1 _8078_ (
  .A(_3497_),
  .ZN(_3498_)
);

NOR3_X1 _8079_ (
  .A1(_3428_),
  .A2(_3394_),
  .A3(_3405_),
  .ZN(_3499_)
);

NAND3_X1 _8080_ (
  .A1(_3499_),
  .A2(_3490_),
  .A3(_3392_),
  .ZN(_3500_)
);

NAND3_X1 _8081_ (
  .A1(_3491_),
  .A2(_3498_),
  .A3(_3500_),
  .ZN(_3501_)
);

NAND2_X1 _8082_ (
  .A1(_3501_),
  .A2(_4497_),
  .ZN(_3502_)
);

INV_X1 _8083_ (
  .A(_4497_),
  .ZN(_3503_)
);

NAND4_X1 _8084_ (
  .A1(_3491_),
  .A2(_3500_),
  .A3(_3498_),
  .A4(_3503_),
  .ZN(_3504_)
);

NAND3_X1 _8085_ (
  .A1(_3502_),
  .A2(_3504_),
  .A3(_2161_),
  .ZN(_3505_)
);

NAND2_X1 _8086_ (
  .A1(_1728_),
  .A2(\s_pipe[7][22] ),
  .ZN(_3506_)
);

NAND2_X1 _8087_ (
  .A1(_3505_),
  .A2(_3506_),
  .ZN(_0598_)
);

NAND2_X1 _8088_ (
  .A1(_4494_),
  .A2(_4497_),
  .ZN(_3507_)
);

OR2_X2 _8089_ (
  .A1(_3507_),
  .A2(_3468_),
  .ZN(_3508_)
);

INV_X1 _8090_ (
  .A(_3508_),
  .ZN(_3509_)
);

NAND2_X1 _8091_ (
  .A1(_3442_),
  .A2(_3509_),
  .ZN(_3510_)
);

INV_X1 _8092_ (
  .A(_4496_),
  .ZN(_3511_)
);

OAI21_X1 _8093_ (
  .A(_3511_),
  .B1(_3503_),
  .B2(_3494_),
  .ZN(_3512_)
);

INV_X1 _8094_ (
  .A(_3512_),
  .ZN(_3513_)
);

OAI21_X1 _8095_ (
  .A(_3513_),
  .B1(_3475_),
  .B2(_3507_),
  .ZN(_3514_)
);

INV_X1 _8096_ (
  .A(_3514_),
  .ZN(_3515_)
);

INV_X1 _8097_ (
  .A(_3404_),
  .ZN(_3516_)
);

NOR2_X1 _8098_ (
  .A1(_3508_),
  .A2(_3436_),
  .ZN(_3517_)
);

NAND2_X1 _8099_ (
  .A1(_3516_),
  .A2(_3517_),
  .ZN(_3518_)
);

INV_X1 _8100_ (
  .A(_4500_),
  .ZN(_3519_)
);

NAND4_X1 _8101_ (
  .A1(_3510_),
  .A2(_3515_),
  .A3(_3518_),
  .A4(_3519_),
  .ZN(_3520_)
);

NAND3_X1 _8102_ (
  .A1(_3510_),
  .A2(_3515_),
  .A3(_3518_),
  .ZN(_3521_)
);

NAND2_X1 _8103_ (
  .A1(_3521_),
  .A2(_4500_),
  .ZN(_3522_)
);

NAND3_X1 _8104_ (
  .A1(_3520_),
  .A2(_3522_),
  .A3(_2161_),
  .ZN(_3523_)
);

NAND2_X1 _8105_ (
  .A1(_1709_),
  .A2(\s_pipe[7][23] ),
  .ZN(_3524_)
);

NAND2_X1 _8106_ (
  .A1(_3523_),
  .A2(_3524_),
  .ZN(_0599_)
);

NAND2_X1 _8107_ (
  .A1(_1709_),
  .A2(\s_pipe[7][24] ),
  .ZN(_3525_)
);

NOR2_X2 _8108_ (
  .A1(_1198_),
  .A2(\d_pipe[6][23] ),
  .ZN(_3526_)
);

NAND2_X4 _8109_ (
  .A1(_1183_),
  .A2(_3526_),
  .ZN(_3527_)
);

NAND2_X4 _8110_ (
  .A1(_3527_),
  .A2(_0651_),
  .ZN(_3528_)
);

INV_X1 _8111_ (
  .A(\s_pipe[6][23] ),
  .ZN(_3529_)
);

NAND2_X4 _8112_ (
  .A1(_3528_),
  .A2(_3529_),
  .ZN(_3530_)
);

NAND3_X2 _8113_ (
  .A1(_3527_),
  .A2(_0651_),
  .A3(\s_pipe[6][23] ),
  .ZN(_3531_)
);

NAND2_X4 _8114_ (
  .A1(_3530_),
  .A2(_3531_),
  .ZN(_3532_)
);

NAND2_X1 _8115_ (
  .A1(_4497_),
  .A2(_4500_),
  .ZN(_3533_)
);

INV_X1 _8116_ (
  .A(_3533_),
  .ZN(_3534_)
);

NAND2_X1 _8117_ (
  .A1(_3495_),
  .A2(_3534_),
  .ZN(_3535_)
);

INV_X1 _8118_ (
  .A(_4499_),
  .ZN(_3536_)
);

OAI21_X1 _8119_ (
  .A(_3536_),
  .B1(_3519_),
  .B2(_3511_),
  .ZN(_3537_)
);

INV_X1 _8120_ (
  .A(_3537_),
  .ZN(_3538_)
);

NAND2_X1 _8121_ (
  .A1(_3535_),
  .A2(_3538_),
  .ZN(_3539_)
);

INV_X1 _8122_ (
  .A(_3539_),
  .ZN(_3540_)
);

NOR2_X2 _8123_ (
  .A1(_3489_),
  .A2(_3533_),
  .ZN(_3541_)
);

NAND2_X1 _8124_ (
  .A1(_3458_),
  .A2(_3541_),
  .ZN(_3542_)
);

NAND2_X2 _8125_ (
  .A1(_3540_),
  .A2(_3542_),
  .ZN(_3543_)
);

NAND2_X1 _8126_ (
  .A1(_3541_),
  .A2(_3451_),
  .ZN(_3544_)
);

AOI21_X2 _8127_ (
  .A(_3544_),
  .B1(_3410_),
  .B2(_3411_),
  .ZN(_3545_)
);

NOR2_X2 _8128_ (
  .A1(_3543_),
  .A2(_3545_),
  .ZN(_3546_)
);

NAND2_X2 _8129_ (
  .A1(_3532_),
  .A2(_3546_),
  .ZN(_3547_)
);

NAND2_X2 _8130_ (
  .A1(_3547_),
  .A2(_1406_),
  .ZN(_3548_)
);

NOR2_X2 _8131_ (
  .A1(_3532_),
  .A2(_3546_),
  .ZN(_3549_)
);

OAI21_X2 _8132_ (
  .A(_3525_),
  .B1(_3548_),
  .B2(_3549_),
  .ZN(_0600_)
);

NAND2_X1 _8133_ (
  .A1(_2349_),
  .A2(\s_pipe[7][7] ),
  .ZN(_3550_)
);

OAI21_X1 _8134_ (
  .A(_3550_),
  .B1(_2291_),
  .B2(_2726_),
  .ZN(_0601_)
);

NAND2_X1 _8135_ (
  .A1(_1899_),
  .A2(\s_pipe[7][8] ),
  .ZN(_3551_)
);

OAI21_X1 _8136_ (
  .A(_3551_),
  .B1(_1548_),
  .B2(_2728_),
  .ZN(_0602_)
);

NAND2_X1 _8137_ (
  .A1(_1546_),
  .A2(\s_pipe[7][9] ),
  .ZN(_3552_)
);

OAI21_X1 _8138_ (
  .A(_3552_),
  .B1(_1548_),
  .B2(_2730_),
  .ZN(_0603_)
);

MUX2_X1 _8139_ (
  .A(\s_pipe[8][11] ),
  .B(\s_pipe[7][10] ),
  .S(_1564_),
  .Z(_0604_)
);

MUX2_X1 _8140_ (
  .A(\s_pipe[8][12] ),
  .B(_0129_),
  .S(_1564_),
  .Z(_0605_)
);

NAND2_X1 _8141_ (
  .A1(_1522_),
  .A2(\s_pipe[8][13] ),
  .ZN(_3553_)
);

OAI21_X1 _8142_ (
  .A(_3553_),
  .B1(_4098_),
  .B2(_2054_),
  .ZN(_0606_)
);

INV_X1 _8143_ (
  .A(_4097_),
  .ZN(_3554_)
);

NAND2_X1 _8144_ (
  .A1(_3554_),
  .A2(_4437_),
  .ZN(_3555_)
);

INV_X2 _8145_ (
  .A(_4437_),
  .ZN(_3556_)
);

NAND2_X1 _8146_ (
  .A1(_3556_),
  .A2(_4097_),
  .ZN(_3557_)
);

NAND3_X1 _8147_ (
  .A1(_3555_),
  .A2(_3557_),
  .A3(_1572_),
  .ZN(_3558_)
);

INV_X1 _8148_ (
  .A(\s_pipe[8][14] ),
  .ZN(_3559_)
);

OAI21_X1 _8149_ (
  .A(_3558_),
  .B1(_1548_),
  .B2(_3559_),
  .ZN(_0607_)
);

NOR2_X1 _8150_ (
  .A1(_2091_),
  .A2(\s_pipe[8][15] ),
  .ZN(_3560_)
);

INV_X1 _8151_ (
  .A(_4436_),
  .ZN(_3561_)
);

INV_X1 _8152_ (
  .A(_4433_),
  .ZN(_3562_)
);

OAI21_X1 _8153_ (
  .A(_3561_),
  .B1(_3556_),
  .B2(_3562_),
  .ZN(_3563_)
);

NAND2_X1 _8154_ (
  .A1(_4437_),
  .A2(_4434_),
  .ZN(_3564_)
);

NOR2_X1 _8155_ (
  .A1(_3564_),
  .A2(_4096_),
  .ZN(_3565_)
);

NOR2_X2 _8156_ (
  .A1(_3563_),
  .A2(_3565_),
  .ZN(_3566_)
);

INV_X1 _8157_ (
  .A(_4440_),
  .ZN(_3567_)
);

XNOR2_X1 _8158_ (
  .A(_3566_),
  .B(_3567_),
  .ZN(_3568_)
);

AOI21_X1 _8159_ (
  .A(_3560_),
  .B1(_3568_),
  .B2(_2265_),
  .ZN(_0608_)
);

NOR2_X1 _8160_ (
  .A1(_1353_),
  .A2(\s_pipe[8][16] ),
  .ZN(_3569_)
);

INV_X1 _8161_ (
  .A(_4439_),
  .ZN(_3570_)
);

OAI21_X2 _8162_ (
  .A(_3570_),
  .B1(_3567_),
  .B2(_3561_),
  .ZN(_3571_)
);

INV_X2 _8163_ (
  .A(_3571_),
  .ZN(_3572_)
);

NAND3_X1 _8164_ (
  .A1(_3554_),
  .A2(_4437_),
  .A3(_4440_),
  .ZN(_3573_)
);

NAND2_X2 _8165_ (
  .A1(_3572_),
  .A2(_3573_),
  .ZN(_3574_)
);

BUF_X4 _8166_ (
  .A(_4443_),
  .Z(_3575_)
);

XNOR2_X1 _8167_ (
  .A(_3574_),
  .B(_3575_),
  .ZN(_3576_)
);

AOI21_X1 _8168_ (
  .A(_3569_),
  .B1(_3576_),
  .B2(_1381_),
  .ZN(_0609_)
);

NOR2_X1 _8169_ (
  .A1(_1371_),
  .A2(\s_pipe[8][17] ),
  .ZN(_3577_)
);

INV_X1 _8170_ (
  .A(_4442_),
  .ZN(_3578_)
);

INV_X1 _8171_ (
  .A(_3575_),
  .ZN(_3579_)
);

OAI21_X1 _8172_ (
  .A(_3578_),
  .B1(_3579_),
  .B2(_3570_),
  .ZN(_3580_)
);

INV_X1 _8173_ (
  .A(_3580_),
  .ZN(_3581_)
);

NAND2_X2 _8174_ (
  .A1(_4440_),
  .A2(_3575_),
  .ZN(_3582_)
);

OAI21_X2 _8175_ (
  .A(_3581_),
  .B1(_3566_),
  .B2(_3582_),
  .ZN(_3583_)
);

BUF_X4 _8176_ (
  .A(_4446_),
  .Z(_3584_)
);

XNOR2_X1 _8177_ (
  .A(_3583_),
  .B(_3584_),
  .ZN(_3585_)
);

AOI21_X1 _8178_ (
  .A(_3577_),
  .B1(_3585_),
  .B2(_1381_),
  .ZN(_0610_)
);

NOR2_X1 _8179_ (
  .A1(_2091_),
  .A2(\s_pipe[8][18] ),
  .ZN(_3586_)
);

NAND2_X2 _8180_ (
  .A1(_3584_),
  .A2(_4442_),
  .ZN(_3587_)
);

INV_X1 _8181_ (
  .A(_4445_),
  .ZN(_3588_)
);

NAND2_X2 _8182_ (
  .A1(_3587_),
  .A2(_3588_),
  .ZN(_3589_)
);

NAND2_X2 _8183_ (
  .A1(_3575_),
  .A2(_3584_),
  .ZN(_3590_)
);

INV_X1 _8184_ (
  .A(_3590_),
  .ZN(_3591_)
);

AOI21_X1 _8185_ (
  .A(_3589_),
  .B1(_3574_),
  .B2(_3591_),
  .ZN(_3592_)
);

INV_X1 _8186_ (
  .A(_4449_),
  .ZN(_3593_)
);

XNOR2_X1 _8187_ (
  .A(_3592_),
  .B(_3593_),
  .ZN(_3594_)
);

AOI21_X1 _8188_ (
  .A(_3586_),
  .B1(_3594_),
  .B2(_1552_),
  .ZN(_0611_)
);

INV_X1 _8189_ (
  .A(_3582_),
  .ZN(_3595_)
);

NAND2_X1 _8190_ (
  .A1(_3584_),
  .A2(_4449_),
  .ZN(_3596_)
);

INV_X1 _8191_ (
  .A(_3596_),
  .ZN(_3597_)
);

NAND2_X1 _8192_ (
  .A1(_3595_),
  .A2(_3597_),
  .ZN(_3598_)
);

OR2_X2 _8193_ (
  .A1(_3566_),
  .A2(_3598_),
  .ZN(_3599_)
);

NAND2_X1 _8194_ (
  .A1(_3580_),
  .A2(_3597_),
  .ZN(_3600_)
);

INV_X1 _8195_ (
  .A(_4448_),
  .ZN(_3601_)
);

OAI21_X1 _8196_ (
  .A(_3601_),
  .B1(_3593_),
  .B2(_3588_),
  .ZN(_3602_)
);

INV_X1 _8197_ (
  .A(_3602_),
  .ZN(_3603_)
);

NAND2_X1 _8198_ (
  .A1(_3600_),
  .A2(_3603_),
  .ZN(_3604_)
);

INV_X1 _8199_ (
  .A(_3604_),
  .ZN(_3605_)
);

NAND2_X1 _8200_ (
  .A1(_3599_),
  .A2(_3605_),
  .ZN(_3606_)
);

NAND2_X1 _8201_ (
  .A1(_3606_),
  .A2(_4452_),
  .ZN(_3607_)
);

INV_X1 _8202_ (
  .A(_4452_),
  .ZN(_3608_)
);

NAND3_X1 _8203_ (
  .A1(_3599_),
  .A2(_3605_),
  .A3(_3608_),
  .ZN(_3609_)
);

NAND3_X1 _8204_ (
  .A1(_3607_),
  .A2(_3609_),
  .A3(_1406_),
  .ZN(_3610_)
);

INV_X1 _8205_ (
  .A(\s_pipe[8][19] ),
  .ZN(_3611_)
);

OAI21_X1 _8206_ (
  .A(_3610_),
  .B1(_1408_),
  .B2(_3611_),
  .ZN(_0612_)
);

NAND2_X2 _8207_ (
  .A1(_4449_),
  .A2(_4452_),
  .ZN(_3612_)
);

NOR2_X2 _8208_ (
  .A1(_3590_),
  .A2(_3612_),
  .ZN(_3613_)
);

NAND2_X1 _8209_ (
  .A1(_3574_),
  .A2(_3613_),
  .ZN(_3614_)
);

INV_X1 _8210_ (
  .A(_4451_),
  .ZN(_3615_)
);

OAI21_X2 _8211_ (
  .A(_3615_),
  .B1(_3608_),
  .B2(_3601_),
  .ZN(_3616_)
);

INV_X1 _8212_ (
  .A(_3616_),
  .ZN(_3617_)
);

INV_X1 _8213_ (
  .A(_3612_),
  .ZN(_3618_)
);

NAND2_X1 _8214_ (
  .A1(_3589_),
  .A2(_3618_),
  .ZN(_3619_)
);

NAND2_X1 _8215_ (
  .A1(_3617_),
  .A2(_3619_),
  .ZN(_3620_)
);

INV_X1 _8216_ (
  .A(_3620_),
  .ZN(_3621_)
);

NAND2_X1 _8217_ (
  .A1(_3614_),
  .A2(_3621_),
  .ZN(_3622_)
);

NAND2_X1 _8218_ (
  .A1(_3622_),
  .A2(_4455_),
  .ZN(_3623_)
);

INV_X1 _8219_ (
  .A(_4455_),
  .ZN(_3624_)
);

NAND3_X1 _8220_ (
  .A1(_3614_),
  .A2(_3624_),
  .A3(_3621_),
  .ZN(_3625_)
);

NAND3_X1 _8221_ (
  .A1(_3623_),
  .A2(_3625_),
  .A3(_1406_),
  .ZN(_3626_)
);

INV_X1 _8222_ (
  .A(\s_pipe[8][20] ),
  .ZN(_3627_)
);

OAI21_X1 _8223_ (
  .A(_3626_),
  .B1(_1634_),
  .B2(_3627_),
  .ZN(_0613_)
);

NAND2_X1 _8224_ (
  .A1(_3563_),
  .A2(_3595_),
  .ZN(_3628_)
);

NAND2_X1 _8225_ (
  .A1(_3628_),
  .A2(_3581_),
  .ZN(_3629_)
);

NAND2_X2 _8226_ (
  .A1(_4452_),
  .A2(_4455_),
  .ZN(_3630_)
);

NOR2_X1 _8227_ (
  .A1(_3596_),
  .A2(_3630_),
  .ZN(_3631_)
);

NAND2_X1 _8228_ (
  .A1(_3629_),
  .A2(_3631_),
  .ZN(_3632_)
);

INV_X1 _8229_ (
  .A(_3630_),
  .ZN(_3633_)
);

NAND2_X1 _8230_ (
  .A1(_3602_),
  .A2(_3633_),
  .ZN(_3634_)
);

INV_X1 _8231_ (
  .A(_4454_),
  .ZN(_3635_)
);

OAI21_X1 _8232_ (
  .A(_3635_),
  .B1(_3624_),
  .B2(_3615_),
  .ZN(_3636_)
);

INV_X1 _8233_ (
  .A(_3636_),
  .ZN(_3637_)
);

NAND2_X1 _8234_ (
  .A1(_3634_),
  .A2(_3637_),
  .ZN(_3638_)
);

INV_X1 _8235_ (
  .A(_3638_),
  .ZN(_3639_)
);

NOR2_X1 _8236_ (
  .A1(_3564_),
  .A2(_3582_),
  .ZN(_3640_)
);

NAND3_X1 _8237_ (
  .A1(_3640_),
  .A2(_3631_),
  .A3(_4100_),
  .ZN(_3641_)
);

NAND3_X1 _8238_ (
  .A1(_3632_),
  .A2(_3639_),
  .A3(_3641_),
  .ZN(_3642_)
);

NAND2_X1 _8239_ (
  .A1(_3642_),
  .A2(_4458_),
  .ZN(_3643_)
);

INV_X1 _8240_ (
  .A(_4458_),
  .ZN(_3644_)
);

NAND4_X1 _8241_ (
  .A1(_3632_),
  .A2(_3641_),
  .A3(_3639_),
  .A4(_3644_),
  .ZN(_3645_)
);

NAND3_X1 _8242_ (
  .A1(_3643_),
  .A2(_3645_),
  .A3(_2349_),
  .ZN(_3646_)
);

NAND2_X1 _8243_ (
  .A1(_1859_),
  .A2(\s_pipe[8][21] ),
  .ZN(_3647_)
);

NAND2_X1 _8244_ (
  .A1(_3646_),
  .A2(_3647_),
  .ZN(_0614_)
);

NAND2_X1 _8245_ (
  .A1(_3571_),
  .A2(_3591_),
  .ZN(_3648_)
);

INV_X1 _8246_ (
  .A(_3589_),
  .ZN(_3649_)
);

NAND2_X1 _8247_ (
  .A1(_3648_),
  .A2(_3649_),
  .ZN(_3650_)
);

NAND2_X1 _8248_ (
  .A1(_4455_),
  .A2(_4458_),
  .ZN(_3651_)
);

NOR2_X1 _8249_ (
  .A1(_3612_),
  .A2(_3651_),
  .ZN(_3652_)
);

NAND2_X1 _8250_ (
  .A1(_3650_),
  .A2(_3652_),
  .ZN(_3653_)
);

INV_X1 _8251_ (
  .A(_3651_),
  .ZN(_3654_)
);

NAND2_X1 _8252_ (
  .A1(_3616_),
  .A2(_3654_),
  .ZN(_3655_)
);

INV_X1 _8253_ (
  .A(_4457_),
  .ZN(_3656_)
);

OAI21_X1 _8254_ (
  .A(_3656_),
  .B1(_3644_),
  .B2(_3635_),
  .ZN(_3657_)
);

INV_X1 _8255_ (
  .A(_3657_),
  .ZN(_3658_)
);

NAND2_X1 _8256_ (
  .A1(_3655_),
  .A2(_3658_),
  .ZN(_3659_)
);

INV_X1 _8257_ (
  .A(_3659_),
  .ZN(_3660_)
);

NOR3_X1 _8258_ (
  .A1(_3590_),
  .A2(_3556_),
  .A3(_3567_),
  .ZN(_3661_)
);

NAND3_X1 _8259_ (
  .A1(_3661_),
  .A2(_3652_),
  .A3(_3554_),
  .ZN(_3662_)
);

NAND3_X1 _8260_ (
  .A1(_3653_),
  .A2(_3660_),
  .A3(_3662_),
  .ZN(_3663_)
);

NAND2_X1 _8261_ (
  .A1(_3663_),
  .A2(_4461_),
  .ZN(_3664_)
);

INV_X1 _8262_ (
  .A(_4461_),
  .ZN(_3665_)
);

NAND4_X1 _8263_ (
  .A1(_3653_),
  .A2(_3662_),
  .A3(_3660_),
  .A4(_3665_),
  .ZN(_3666_)
);

NAND3_X1 _8264_ (
  .A1(_3664_),
  .A2(_3666_),
  .A3(_1447_),
  .ZN(_3667_)
);

NAND2_X1 _8265_ (
  .A1(_1859_),
  .A2(\s_pipe[8][22] ),
  .ZN(_3668_)
);

NAND2_X1 _8266_ (
  .A1(_3667_),
  .A2(_3668_),
  .ZN(_0615_)
);

NAND2_X1 _8267_ (
  .A1(_4458_),
  .A2(_4461_),
  .ZN(_3669_)
);

OR2_X2 _8268_ (
  .A1(_3669_),
  .A2(_3630_),
  .ZN(_3670_)
);

INV_X1 _8269_ (
  .A(_3670_),
  .ZN(_3671_)
);

NAND2_X1 _8270_ (
  .A1(_3604_),
  .A2(_3671_),
  .ZN(_3672_)
);

INV_X1 _8271_ (
  .A(_4460_),
  .ZN(_3673_)
);

OAI21_X1 _8272_ (
  .A(_3673_),
  .B1(_3665_),
  .B2(_3656_),
  .ZN(_3674_)
);

INV_X1 _8273_ (
  .A(_3674_),
  .ZN(_3675_)
);

OAI21_X1 _8274_ (
  .A(_3675_),
  .B1(_3637_),
  .B2(_3669_),
  .ZN(_3676_)
);

INV_X1 _8275_ (
  .A(_3676_),
  .ZN(_3677_)
);

INV_X1 _8276_ (
  .A(_3566_),
  .ZN(_3678_)
);

NOR2_X2 _8277_ (
  .A1(_3670_),
  .A2(_3598_),
  .ZN(_3679_)
);

NAND2_X1 _8278_ (
  .A1(_3678_),
  .A2(_3679_),
  .ZN(_3680_)
);

INV_X1 _8279_ (
  .A(_4464_),
  .ZN(_3681_)
);

NAND4_X1 _8280_ (
  .A1(_3672_),
  .A2(_3677_),
  .A3(_3680_),
  .A4(_3681_),
  .ZN(_3682_)
);

NAND3_X1 _8281_ (
  .A1(_3672_),
  .A2(_3677_),
  .A3(_3680_),
  .ZN(_3683_)
);

NAND2_X1 _8282_ (
  .A1(_3683_),
  .A2(_4464_),
  .ZN(_3684_)
);

NAND3_X1 _8283_ (
  .A1(_3682_),
  .A2(_3684_),
  .A3(_2001_),
  .ZN(_3685_)
);

NAND2_X1 _8284_ (
  .A1(_1728_),
  .A2(\s_pipe[8][23] ),
  .ZN(_3686_)
);

NAND2_X1 _8285_ (
  .A1(_3685_),
  .A2(_3686_),
  .ZN(_0616_)
);

NAND2_X1 _8286_ (
  .A1(_1522_),
  .A2(\s_pipe[8][24] ),
  .ZN(_3687_)
);

NOR2_X1 _8287_ (
  .A1(_1138_),
  .A2(\d_pipe[7][23] ),
  .ZN(_3688_)
);

NAND2_X2 _8288_ (
  .A1(_1122_),
  .A2(_3688_),
  .ZN(_3689_)
);

NAND2_X1 _8289_ (
  .A1(_3689_),
  .A2(_0648_),
  .ZN(_3690_)
);

INV_X1 _8290_ (
  .A(\s_pipe[7][23] ),
  .ZN(_3691_)
);

NAND2_X1 _8291_ (
  .A1(_3690_),
  .A2(_3691_),
  .ZN(_3692_)
);

NAND3_X1 _8292_ (
  .A1(_3689_),
  .A2(_0648_),
  .A3(\s_pipe[7][23] ),
  .ZN(_3693_)
);

NAND2_X2 _8293_ (
  .A1(_3692_),
  .A2(_3693_),
  .ZN(_3694_)
);

NAND2_X1 _8294_ (
  .A1(_4461_),
  .A2(_4464_),
  .ZN(_3695_)
);

INV_X1 _8295_ (
  .A(_3695_),
  .ZN(_3696_)
);

NAND2_X1 _8296_ (
  .A1(_3657_),
  .A2(_3696_),
  .ZN(_3697_)
);

INV_X1 _8297_ (
  .A(_4463_),
  .ZN(_3698_)
);

OAI21_X1 _8298_ (
  .A(_3698_),
  .B1(_3681_),
  .B2(_3673_),
  .ZN(_3699_)
);

INV_X1 _8299_ (
  .A(_3699_),
  .ZN(_3700_)
);

NAND2_X1 _8300_ (
  .A1(_3697_),
  .A2(_3700_),
  .ZN(_3701_)
);

INV_X1 _8301_ (
  .A(_3701_),
  .ZN(_3702_)
);

NOR2_X2 _8302_ (
  .A1(_3651_),
  .A2(_3695_),
  .ZN(_3703_)
);

NAND2_X1 _8303_ (
  .A1(_3620_),
  .A2(_3703_),
  .ZN(_3704_)
);

NAND2_X1 _8304_ (
  .A1(_3702_),
  .A2(_3704_),
  .ZN(_3705_)
);

NAND2_X1 _8305_ (
  .A1(_3703_),
  .A2(_3613_),
  .ZN(_3706_)
);

AOI21_X2 _8306_ (
  .A(_3706_),
  .B1(_3572_),
  .B2(_3573_),
  .ZN(_3707_)
);

NOR2_X1 _8307_ (
  .A1(_3705_),
  .A2(_3707_),
  .ZN(_3708_)
);

NAND2_X1 _8308_ (
  .A1(_3694_),
  .A2(_3708_),
  .ZN(_3709_)
);

NAND2_X1 _8309_ (
  .A1(_3709_),
  .A2(_1406_),
  .ZN(_3710_)
);

NOR2_X1 _8310_ (
  .A1(_3694_),
  .A2(_3708_),
  .ZN(_3711_)
);

OAI21_X2 _8311_ (
  .A(_3687_),
  .B1(_3710_),
  .B2(_3711_),
  .ZN(_0617_)
);

FA_X1 _8312_ (
  .A(_4042_),
  .B(_4043_),
  .CI(_4044_),
  .CO(_4045_),
  .S(_4046_)
);

FA_X1 _8313_ (
  .A(_4049_),
  .B(_4050_),
  .CI(_4051_),
  .CO(_4052_),
  .S(_4053_)
);

FA_X1 _8314_ (
  .A(_4056_),
  .B(_4057_),
  .CI(_4058_),
  .CO(_4059_),
  .S(_4060_)
);

FA_X1 _8315_ (
  .A(_4063_),
  .B(d[1]),
  .CI(_4064_),
  .CO(_4065_),
  .S(_0143_)
);

FA_X1 _8316_ (
  .A(_4066_),
  .B(_4067_),
  .CI(_4068_),
  .CO(_4069_),
  .S(_4070_)
);

FA_X1 _8317_ (
  .A(_4073_),
  .B(_4074_),
  .CI(_4075_),
  .CO(_4076_),
  .S(_4077_)
);

FA_X1 _8318_ (
  .A(_4080_),
  .B(_4081_),
  .CI(_4082_),
  .CO(_4083_),
  .S(_4084_)
);

FA_X1 _8319_ (
  .A(_4087_),
  .B(_4088_),
  .CI(_4089_),
  .CO(_4090_),
  .S(_4091_)
);

FA_X1 _8320_ (
  .A(_4094_),
  .B(_4095_),
  .CI(_4096_),
  .CO(_4097_),
  .S(_4098_)
);

FA_X1 _8321_ (
  .A(_4101_),
  .B(_4102_),
  .CI(_4103_),
  .CO(_4104_),
  .S(_4105_)
);

FA_X1 _8322_ (
  .A(_4108_),
  .B(_4109_),
  .CI(_4110_),
  .CO(_4111_),
  .S(_4112_)
);

FA_X1 _8323_ (
  .A(_4115_),
  .B(_4116_),
  .CI(_4117_),
  .CO(_4118_),
  .S(_4119_)
);

HA_X1 _8324_ (
  .A(_4122_),
  .B(d[0]),
  .CO(_4064_),
  .S(_4123_)
);

HA_X1 _8335_ (
  .A(_4144_),
  .B(_4145_),
  .CO(_4146_),
  .S(_4147_)
);

HA_X1 _8336_ (
  .A(\s_pipe[2][12] ),
  .B(_4048_),
  .CO(_4148_),
  .S(_4149_)
);

HA_X1 _8337_ (
  .A(\s_pipe[2][13] ),
  .B(_4150_),
  .CO(_4151_),
  .S(_4152_)
);

HA_X1 _8338_ (
  .A(\s_pipe[2][14] ),
  .B(_4153_),
  .CO(_4154_),
  .S(_4155_)
);

HA_X1 _8339_ (
  .A(\s_pipe[2][15] ),
  .B(_4156_),
  .CO(_4157_),
  .S(_4158_)
);

HA_X1 _8340_ (
  .A(\s_pipe[2][16] ),
  .B(_4159_),
  .CO(_4160_),
  .S(_4161_)
);

HA_X1 _8341_ (
  .A(\s_pipe[2][17] ),
  .B(_4162_),
  .CO(_4163_),
  .S(_4164_)
);

HA_X1 _8342_ (
  .A(\s_pipe[2][18] ),
  .B(_4165_),
  .CO(_4166_),
  .S(_4167_)
);

HA_X1 _8343_ (
  .A(\s_pipe[2][19] ),
  .B(_4168_),
  .CO(_4169_),
  .S(_4170_)
);

HA_X1 _8344_ (
  .A(\s_pipe[2][20] ),
  .B(_4171_),
  .CO(_4172_),
  .S(_4173_)
);

HA_X1 _8345_ (
  .A(\s_pipe[2][21] ),
  .B(_4174_),
  .CO(_4175_),
  .S(_4176_)
);

HA_X1 _8346_ (
  .A(\s_pipe[2][22] ),
  .B(_4177_),
  .CO(_4178_),
  .S(_4179_)
);

HA_X1 _8347_ (
  .A(\d_pipe[3][12] ),
  .B(\s_pipe[3][11] ),
  .CO(_4054_),
  .S(_0125_)
);

HA_X1 _8348_ (
  .A(_4180_),
  .B(_4181_),
  .CO(_4182_),
  .S(_4183_)
);

HA_X1 _8349_ (
  .A(\s_pipe[3][12] ),
  .B(_4055_),
  .CO(_4184_),
  .S(_4185_)
);

HA_X1 _8350_ (
  .A(\s_pipe[3][13] ),
  .B(_4186_),
  .CO(_4187_),
  .S(_4188_)
);

HA_X1 _8351_ (
  .A(\s_pipe[3][14] ),
  .B(_4189_),
  .CO(_4190_),
  .S(_4191_)
);

HA_X1 _8352_ (
  .A(\s_pipe[3][15] ),
  .B(_4192_),
  .CO(_4193_),
  .S(_4194_)
);

HA_X1 _8353_ (
  .A(\s_pipe[3][16] ),
  .B(_4195_),
  .CO(_4196_),
  .S(_4197_)
);

HA_X1 _8354_ (
  .A(\s_pipe[3][17] ),
  .B(_4198_),
  .CO(_4199_),
  .S(_4200_)
);

HA_X1 _8355_ (
  .A(\s_pipe[3][18] ),
  .B(_4201_),
  .CO(_4202_),
  .S(_4203_)
);

HA_X1 _8356_ (
  .A(\s_pipe[3][19] ),
  .B(_4204_),
  .CO(_4205_),
  .S(_4206_)
);

HA_X1 _8357_ (
  .A(\s_pipe[3][20] ),
  .B(_4207_),
  .CO(_4208_),
  .S(_4209_)
);

HA_X1 _8358_ (
  .A(\s_pipe[3][21] ),
  .B(_4210_),
  .CO(_4211_),
  .S(_4212_)
);

HA_X1 _8359_ (
  .A(\s_pipe[3][22] ),
  .B(_4213_),
  .CO(_4214_),
  .S(_4215_)
);

HA_X1 _8360_ (
  .A(\d_pipe[1][12] ),
  .B(\s_pipe[1][11] ),
  .CO(_4062_),
  .S(_0123_)
);

HA_X1 _8361_ (
  .A(_4216_),
  .B(_4217_),
  .CO(_4218_),
  .S(_4219_)
);

HA_X1 _8362_ (
  .A(\s_pipe[1][12] ),
  .B(_4061_),
  .CO(_4220_),
  .S(_4221_)
);

HA_X1 _8363_ (
  .A(\s_pipe[1][13] ),
  .B(_4222_),
  .CO(_4223_),
  .S(_4224_)
);

HA_X1 _8364_ (
  .A(\s_pipe[1][14] ),
  .B(_4225_),
  .CO(_4226_),
  .S(_4227_)
);

HA_X1 _8365_ (
  .A(\s_pipe[1][15] ),
  .B(_4228_),
  .CO(_4229_),
  .S(_4230_)
);

HA_X1 _8366_ (
  .A(\s_pipe[1][16] ),
  .B(_4231_),
  .CO(_4232_),
  .S(_4233_)
);

HA_X1 _8367_ (
  .A(\s_pipe[1][17] ),
  .B(_4234_),
  .CO(_4235_),
  .S(_4236_)
);

HA_X1 _8368_ (
  .A(\s_pipe[1][18] ),
  .B(_4237_),
  .CO(_4238_),
  .S(_4239_)
);

HA_X1 _8369_ (
  .A(\s_pipe[1][19] ),
  .B(_4240_),
  .CO(_4241_),
  .S(_4242_)
);

HA_X1 _8370_ (
  .A(\s_pipe[1][20] ),
  .B(_4243_),
  .CO(_4244_),
  .S(_4245_)
);

HA_X1 _8371_ (
  .A(\s_pipe[1][21] ),
  .B(_4246_),
  .CO(_4247_),
  .S(_4248_)
);

HA_X1 _8372_ (
  .A(\s_pipe[1][22] ),
  .B(_4249_),
  .CO(_4250_),
  .S(_4251_)
);

HA_X1 _8373_ (
  .A(z[12]),
  .B(_4252_),
  .CO(_4253_),
  .S(_4254_)
);

HA_X1 _8374_ (
  .A(z[13]),
  .B(_4255_),
  .CO(_4256_),
  .S(_4257_)
);

HA_X1 _8375_ (
  .A(z[14]),
  .B(_4258_),
  .CO(_4259_),
  .S(_4260_)
);

HA_X1 _8376_ (
  .A(z[15]),
  .B(_4261_),
  .CO(_4262_),
  .S(_4263_)
);

HA_X1 _8377_ (
  .A(z[16]),
  .B(_4264_),
  .CO(_4265_),
  .S(_4266_)
);

HA_X1 _8378_ (
  .A(z[17]),
  .B(_4267_),
  .CO(_4268_),
  .S(_4269_)
);

HA_X1 _8379_ (
  .A(z[18]),
  .B(_4270_),
  .CO(_4271_),
  .S(_4272_)
);

HA_X1 _8380_ (
  .A(z[19]),
  .B(_4273_),
  .CO(_4274_),
  .S(_4275_)
);

HA_X1 _8381_ (
  .A(z[20]),
  .B(_4276_),
  .CO(_4277_),
  .S(_4278_)
);

HA_X1 _8382_ (
  .A(z[21]),
  .B(_4279_),
  .CO(_4280_),
  .S(_4281_)
);

HA_X1 _8383_ (
  .A(z[22]),
  .B(_4282_),
  .CO(_4283_),
  .S(_4284_)
);

HA_X1 _8384_ (
  .A(\d_pipe[11][12] ),
  .B(\s_pipe[11][11] ),
  .CO(_4072_),
  .S(_0142_)
);

HA_X1 _8385_ (
  .A(_4285_),
  .B(_4286_),
  .CO(_4287_),
  .S(_4288_)
);

HA_X1 _8387_ (
  .A(\s_pipe[11][13] ),
  .B(_4291_),
  .CO(_4292_),
  .S(_4293_)
);

HA_X1 _8388_ (
  .A(\s_pipe[11][14] ),
  .B(_4294_),
  .CO(_4295_),
  .S(_4296_)
);

HA_X1 _8389_ (
  .A(\s_pipe[11][15] ),
  .B(_4297_),
  .CO(_4298_),
  .S(_4299_)
);

HA_X1 _8390_ (
  .A(\s_pipe[11][16] ),
  .B(_4300_),
  .CO(_4301_),
  .S(_4302_)
);

HA_X1 _8391_ (
  .A(\s_pipe[11][17] ),
  .B(_4303_),
  .CO(_4304_),
  .S(_4305_)
);

HA_X1 _8392_ (
  .A(\s_pipe[11][18] ),
  .B(_4306_),
  .CO(_4307_),
  .S(_4308_)
);

HA_X1 _8393_ (
  .A(\s_pipe[11][19] ),
  .B(_4309_),
  .CO(_4310_),
  .S(_4311_)
);

HA_X1 _8394_ (
  .A(\s_pipe[11][20] ),
  .B(_4312_),
  .CO(_4313_),
  .S(_4314_)
);

HA_X1 _8395_ (
  .A(\s_pipe[11][21] ),
  .B(_4315_),
  .CO(_4316_),
  .S(_4317_)
);

HA_X1 _8396_ (
  .A(\s_pipe[11][22] ),
  .B(_4318_),
  .CO(_4319_),
  .S(_4320_)
);

HA_X1 _8397_ (
  .A(\d_pipe[10][12] ),
  .B(\s_pipe[10][11] ),
  .CO(_4079_),
  .S(_0141_)
);

HA_X1 _8398_ (
  .A(_4321_),
  .B(_4322_),
  .CO(_4323_),
  .S(_4324_)
);

HA_X1 _8399_ (
  .A(\s_pipe[10][12] ),
  .B(_4078_),
  .CO(_4325_),
  .S(_4326_)
);

HA_X1 _8400_ (
  .A(\s_pipe[10][13] ),
  .B(_4327_),
  .CO(_4328_),
  .S(_4329_)
);

HA_X1 _8401_ (
  .A(\s_pipe[10][14] ),
  .B(_4330_),
  .CO(_4331_),
  .S(_4332_)
);

HA_X1 _8402_ (
  .A(\s_pipe[10][15] ),
  .B(_4333_),
  .CO(_4334_),
  .S(_4335_)
);

HA_X1 _8403_ (
  .A(\s_pipe[10][16] ),
  .B(_4336_),
  .CO(_4337_),
  .S(_4338_)
);

HA_X1 _8404_ (
  .A(\s_pipe[10][17] ),
  .B(_4339_),
  .CO(_4340_),
  .S(_4341_)
);

HA_X1 _8405_ (
  .A(\s_pipe[10][18] ),
  .B(_4342_),
  .CO(_4343_),
  .S(_4344_)
);

HA_X1 _8406_ (
  .A(\s_pipe[10][19] ),
  .B(_4345_),
  .CO(_4346_),
  .S(_4347_)
);

HA_X1 _8407_ (
  .A(\s_pipe[10][20] ),
  .B(_4348_),
  .CO(_4349_),
  .S(_4350_)
);

HA_X1 _8408_ (
  .A(\s_pipe[10][21] ),
  .B(_4351_),
  .CO(_4352_),
  .S(_4353_)
);

HA_X1 _8409_ (
  .A(\s_pipe[10][22] ),
  .B(_4354_),
  .CO(_4355_),
  .S(_4356_)
);

HA_X1 _8410_ (
  .A(\d_pipe[9][12] ),
  .B(\s_pipe[9][11] ),
  .CO(_4086_),
  .S(_0140_)
);

HA_X1 _8411_ (
  .A(_4357_),
  .B(_4358_),
  .CO(_4359_),
  .S(_4360_)
);

HA_X1 _8412_ (
  .A(\s_pipe[9][12] ),
  .B(_4085_),
  .CO(_4361_),
  .S(_4362_)
);

HA_X1 _8413_ (
  .A(\s_pipe[9][13] ),
  .B(_4363_),
  .CO(_4364_),
  .S(_4365_)
);

HA_X1 _8414_ (
  .A(\s_pipe[9][14] ),
  .B(_4366_),
  .CO(_4367_),
  .S(_4368_)
);

HA_X1 _8415_ (
  .A(_4369_),
  .B(_0134_),
  .CO(_4370_),
  .S(_4371_)
);

HA_X1 _8416_ (
  .A(_0135_),
  .B(_4372_),
  .CO(_4373_),
  .S(_4374_)
);

HA_X1 _8417_ (
  .A(_0136_),
  .B(_4375_),
  .CO(_4376_),
  .S(_4377_)
);

HA_X1 _8418_ (
  .A(_0137_),
  .B(_4378_),
  .CO(_4379_),
  .S(_4380_)
);

HA_X1 _8419_ (
  .A(_0138_),
  .B(_4381_),
  .CO(_4382_),
  .S(_4383_)
);

HA_X1 _8420_ (
  .A(_0139_),
  .B(_4384_),
  .CO(_4385_),
  .S(_4386_)
);

HA_X1 _8421_ (
  .A(_0131_),
  .B(_4387_),
  .CO(_4388_),
  .S(_4389_)
);

HA_X1 _8422_ (
  .A(_0132_),
  .B(_4390_),
  .CO(_4391_),
  .S(_4392_)
);

HA_X1 _8423_ (
  .A(\d_pipe[8][12] ),
  .B(\s_pipe[8][11] ),
  .CO(_4093_),
  .S(_0130_)
);

HA_X1 _8424_ (
  .A(_4393_),
  .B(_4394_),
  .CO(_4395_),
  .S(_4396_)
);

HA_X1 _8425_ (
  .A(\s_pipe[8][12] ),
  .B(_4092_),
  .CO(_4397_),
  .S(_4398_)
);

HA_X1 _8426_ (
  .A(\s_pipe[8][13] ),
  .B(_4399_),
  .CO(_4400_),
  .S(_4401_)
);

HA_X1 _8427_ (
  .A(\s_pipe[8][14] ),
  .B(_4402_),
  .CO(_4403_),
  .S(_4404_)
);

HA_X1 _8428_ (
  .A(\s_pipe[8][15] ),
  .B(_4405_),
  .CO(_4406_),
  .S(_4407_)
);

HA_X1 _8429_ (
  .A(\s_pipe[8][16] ),
  .B(_4408_),
  .CO(_4409_),
  .S(_4410_)
);

HA_X1 _8430_ (
  .A(\s_pipe[8][17] ),
  .B(_4411_),
  .CO(_4412_),
  .S(_4413_)
);

HA_X1 _8431_ (
  .A(\s_pipe[8][18] ),
  .B(_4414_),
  .CO(_4415_),
  .S(_4416_)
);

HA_X1 _8432_ (
  .A(\s_pipe[8][19] ),
  .B(_4417_),
  .CO(_4418_),
  .S(_4419_)
);

HA_X1 _8433_ (
  .A(\s_pipe[8][20] ),
  .B(_4420_),
  .CO(_4421_),
  .S(_4422_)
);

HA_X1 _8434_ (
  .A(\s_pipe[8][21] ),
  .B(_4423_),
  .CO(_4424_),
  .S(_4425_)
);

HA_X1 _8435_ (
  .A(\s_pipe[8][22] ),
  .B(_4426_),
  .CO(_4427_),
  .S(_4428_)
);

HA_X1 _8436_ (
  .A(\d_pipe[7][12] ),
  .B(\s_pipe[7][11] ),
  .CO(_4100_),
  .S(_0129_)
);

HA_X1 _8437_ (
  .A(_4429_),
  .B(_4430_),
  .CO(_4431_),
  .S(_4432_)
);

HA_X1 _8438_ (
  .A(\s_pipe[7][12] ),
  .B(_4099_),
  .CO(_4433_),
  .S(_4434_)
);

HA_X1 _8439_ (
  .A(\s_pipe[7][13] ),
  .B(_4435_),
  .CO(_4436_),
  .S(_4437_)
);

HA_X1 _8440_ (
  .A(\s_pipe[7][14] ),
  .B(_4438_),
  .CO(_4439_),
  .S(_4440_)
);

HA_X1 _8441_ (
  .A(\s_pipe[7][15] ),
  .B(_4441_),
  .CO(_4442_),
  .S(_4443_)
);

HA_X1 _8442_ (
  .A(\s_pipe[7][16] ),
  .B(_4444_),
  .CO(_4445_),
  .S(_4446_)
);

HA_X1 _8443_ (
  .A(\s_pipe[7][17] ),
  .B(_4447_),
  .CO(_4448_),
  .S(_4449_)
);

HA_X1 _8444_ (
  .A(\s_pipe[7][18] ),
  .B(_4450_),
  .CO(_4451_),
  .S(_4452_)
);

HA_X1 _8445_ (
  .A(\s_pipe[7][19] ),
  .B(_4453_),
  .CO(_4454_),
  .S(_4455_)
);

HA_X1 _8446_ (
  .A(\s_pipe[7][20] ),
  .B(_4456_),
  .CO(_4457_),
  .S(_4458_)
);

HA_X1 _8447_ (
  .A(\s_pipe[7][21] ),
  .B(_4459_),
  .CO(_4460_),
  .S(_4461_)
);

HA_X1 _8448_ (
  .A(\s_pipe[7][22] ),
  .B(_4462_),
  .CO(_4463_),
  .S(_4464_)
);

HA_X1 _8449_ (
  .A(\d_pipe[6][12] ),
  .B(\s_pipe[6][11] ),
  .CO(_4107_),
  .S(_0128_)
);

HA_X1 _8450_ (
  .A(_4465_),
  .B(_4466_),
  .CO(_4467_),
  .S(_4468_)
);

HA_X1 _8451_ (
  .A(\s_pipe[6][12] ),
  .B(_4106_),
  .CO(_4469_),
  .S(_4470_)
);

HA_X1 _8452_ (
  .A(\s_pipe[6][13] ),
  .B(_4471_),
  .CO(_4472_),
  .S(_4473_)
);

HA_X1 _8453_ (
  .A(\s_pipe[6][14] ),
  .B(_4474_),
  .CO(_4475_),
  .S(_4476_)
);

HA_X1 _8454_ (
  .A(\s_pipe[6][15] ),
  .B(_4477_),
  .CO(_4478_),
  .S(_4479_)
);

HA_X1 _8455_ (
  .A(\s_pipe[6][16] ),
  .B(_4480_),
  .CO(_4481_),
  .S(_4482_)
);

HA_X1 _8456_ (
  .A(\s_pipe[6][17] ),
  .B(_4483_),
  .CO(_4484_),
  .S(_4485_)
);

HA_X1 _8457_ (
  .A(\s_pipe[6][18] ),
  .B(_4486_),
  .CO(_4487_),
  .S(_4488_)
);

HA_X1 _8458_ (
  .A(\s_pipe[6][19] ),
  .B(_4489_),
  .CO(_4490_),
  .S(_4491_)
);

HA_X1 _8459_ (
  .A(\s_pipe[6][20] ),
  .B(_4492_),
  .CO(_4493_),
  .S(_4494_)
);

HA_X1 _8460_ (
  .A(\s_pipe[6][21] ),
  .B(_4495_),
  .CO(_4496_),
  .S(_4497_)
);

HA_X1 _8461_ (
  .A(\s_pipe[6][22] ),
  .B(_4498_),
  .CO(_4499_),
  .S(_4500_)
);

HA_X1 _8462_ (
  .A(\d_pipe[5][12] ),
  .B(\s_pipe[5][11] ),
  .CO(_4114_),
  .S(_0127_)
);

HA_X1 _8463_ (
  .A(_4501_),
  .B(_4502_),
  .CO(_4503_),
  .S(_4504_)
);

HA_X1 _8464_ (
  .A(\s_pipe[5][12] ),
  .B(_4113_),
  .CO(_4505_),
  .S(_4506_)
);

HA_X1 _8465_ (
  .A(\s_pipe[5][13] ),
  .B(_4507_),
  .CO(_4508_),
  .S(_4509_)
);

HA_X1 _8466_ (
  .A(\s_pipe[5][14] ),
  .B(_4510_),
  .CO(_4511_),
  .S(_4512_)
);

HA_X1 _8467_ (
  .A(\s_pipe[5][15] ),
  .B(_4513_),
  .CO(_4514_),
  .S(_4515_)
);

HA_X1 _8468_ (
  .A(\s_pipe[5][16] ),
  .B(_4516_),
  .CO(_4517_),
  .S(_4518_)
);

HA_X1 _8469_ (
  .A(\s_pipe[5][17] ),
  .B(_4519_),
  .CO(_4520_),
  .S(_4521_)
);

HA_X1 _8470_ (
  .A(\s_pipe[5][18] ),
  .B(_4522_),
  .CO(_4523_),
  .S(_4524_)
);

HA_X1 _8471_ (
  .A(\s_pipe[5][19] ),
  .B(_4525_),
  .CO(_4526_),
  .S(_4527_)
);

HA_X1 _8472_ (
  .A(\s_pipe[5][20] ),
  .B(_4528_),
  .CO(_4529_),
  .S(_4530_)
);

HA_X1 _8473_ (
  .A(\s_pipe[5][21] ),
  .B(_4531_),
  .CO(_4532_),
  .S(_4533_)
);

HA_X1 _8474_ (
  .A(\s_pipe[5][22] ),
  .B(_4534_),
  .CO(_4535_),
  .S(_4536_)
);

HA_X1 _8475_ (
  .A(\d_pipe[4][12] ),
  .B(\s_pipe[4][11] ),
  .CO(_4121_),
  .S(_0126_)
);

HA_X1 _8476_ (
  .A(_4537_),
  .B(_4538_),
  .CO(_4539_),
  .S(_4540_)
);

HA_X1 _8477_ (
  .A(\s_pipe[4][12] ),
  .B(_4120_),
  .CO(_4541_),
  .S(_4542_)
);

HA_X1 _8478_ (
  .A(\s_pipe[4][13] ),
  .B(_4543_),
  .CO(_4544_),
  .S(_4545_)
);

HA_X1 _8479_ (
  .A(\s_pipe[4][14] ),
  .B(_4546_),
  .CO(_4547_),
  .S(_4548_)
);

HA_X1 _8480_ (
  .A(\s_pipe[4][15] ),
  .B(_4549_),
  .CO(_4550_),
  .S(_4551_)
);

HA_X1 _8481_ (
  .A(\s_pipe[4][16] ),
  .B(_4552_),
  .CO(_4553_),
  .S(_4554_)
);

HA_X1 _8482_ (
  .A(\s_pipe[4][17] ),
  .B(_4555_),
  .CO(_4556_),
  .S(_4557_)
);

HA_X1 _8483_ (
  .A(\s_pipe[4][18] ),
  .B(_4558_),
  .CO(_4559_),
  .S(_4560_)
);

HA_X1 _8484_ (
  .A(\s_pipe[4][19] ),
  .B(_4561_),
  .CO(_4562_),
  .S(_4563_)
);

HA_X1 _8485_ (
  .A(\s_pipe[4][20] ),
  .B(_4564_),
  .CO(_4565_),
  .S(_4566_)
);

HA_X1 _8486_ (
  .A(\s_pipe[4][21] ),
  .B(_4567_),
  .CO(_4568_),
  .S(_4569_)
);

HA_X1 _8487_ (
  .A(\s_pipe[4][22] ),
  .B(_4570_),
  .CO(_4571_),
  .S(_4572_)
);

HA_X1 _8488_ (
  .A(\d_pipe[2][12] ),
  .B(\s_pipe[2][11] ),
  .CO(_4047_),
  .S(_0124_)
);

DFF_X1 _8500_ (
  .D(_0321_),
  .CK(clk),
  .Q(_3714_),
  .QN(_4358_)
);

DFF_X1 _8501_ (
  .D(_0322_),
  .CK(clk),
  .Q(_3715_),
  .QN(_0031_)
);

DFF_X1 _8502_ (
  .D(_0323_),
  .CK(clk),
  .Q(_3716_),
  .QN(_0032_)
);

DFF_X1 _8503_ (
  .D(_0324_),
  .CK(clk),
  .Q(_3717_),
  .QN(_0033_)
);

DFF_X1 _8504_ (
  .D(_0325_),
  .CK(clk),
  .Q(_3718_),
  .QN(_0034_)
);

DFF_X1 _8505_ (
  .D(_0326_),
  .CK(clk),
  .Q(_3719_),
  .QN(_0035_)
);

DFF_X1 _8506_ (
  .D(_0327_),
  .CK(clk),
  .Q(_3720_),
  .QN(_0036_)
);

DFF_X1 _8507_ (
  .D(_0328_),
  .CK(clk),
  .Q(_3721_),
  .QN(_0037_)
);

DFF_X1 _8508_ (
  .D(_0329_),
  .CK(clk),
  .Q(_3722_),
  .QN(_0038_)
);

DFF_X1 _8509_ (
  .D(_0330_),
  .CK(clk),
  .Q(_3712_),
  .QN(_0039_)
);

DFF_X1 _8510_ (
  .D(_0331_),
  .CK(clk),
  .Q(_3713_),
  .QN(_0040_)
);

DFF_X1 _8511_ (
  .D(_0454_),
  .CK(clk),
  .Q(_0134_),
  .QN(_3875_)
);

DFF_X1 _8512_ (
  .D(_0455_),
  .CK(clk),
  .Q(_0135_),
  .QN(_3874_)
);

DFF_X1 _8513_ (
  .D(_0456_),
  .CK(clk),
  .Q(_0136_),
  .QN(_3873_)
);

DFF_X1 _8514_ (
  .D(_0457_),
  .CK(clk),
  .Q(_0137_),
  .QN(_3872_)
);

DFF_X1 _8515_ (
  .D(_0458_),
  .CK(clk),
  .Q(_0138_),
  .QN(_3871_)
);

DFF_X1 _8516_ (
  .D(_0459_),
  .CK(clk),
  .Q(_0139_),
  .QN(_3870_)
);

DFF_X1 _8517_ (
  .D(_0460_),
  .CK(clk),
  .Q(_0131_),
  .QN(_3869_)
);

DFF_X1 _8518_ (
  .D(_0461_),
  .CK(clk),
  .Q(_0132_),
  .QN(_3868_)
);

DFF_X1 _8519_ (
  .D(_0462_),
  .CK(clk),
  .Q(_0133_),
  .QN(_3867_)
);

DFF_X1 _8520_ (
  .D(_0463_),
  .CK(clk),
  .Q(_0000_),
  .QN(_0119_)
);

DFF_X1 _8521_ (
  .D(_0554_),
  .CK(clk),
  .Q(_0618_),
  .QN(_3782_)
);

DFF_X1 _8522_ (
  .D(_0555_),
  .CK(clk),
  .Q(_0619_),
  .QN(_3781_)
);

DFF_X1 _8523_ (
  .D(_0556_),
  .CK(clk),
  .Q(_0620_),
  .QN(_3780_)
);

DFF_X1 _8524_ (
  .D(_0557_),
  .CK(clk),
  .Q(_0621_),
  .QN(_3779_)
);

DFF_X1 _8525_ (
  .D(_0558_),
  .CK(clk),
  .Q(_0622_),
  .QN(_3778_)
);

DFF_X1 _8526_ (
  .D(_0559_),
  .CK(clk),
  .Q(_0623_),
  .QN(_3777_)
);

DFF_X1 _8527_ (
  .D(_0560_),
  .CK(clk),
  .Q(_0624_),
  .QN(_3776_)
);

DFF_X1 _8528_ (
  .D(_0561_),
  .CK(clk),
  .Q(_0625_),
  .QN(_3775_)
);

DFF_X1 \d_pipe[10][12]$_DFFE_PP_  (
  .D(_0332_),
  .CK(clk),
  .Q(\d_pipe[10][12] ),
  .QN(_4321_)
);

DFF_X1 \d_pipe[10][13]$_DFFE_PP_  (
  .D(_0333_),
  .CK(clk),
  .Q(\d_pipe[10][13] ),
  .QN(_4322_)
);

DFF_X1 \d_pipe[10][14]$_DFFE_PP_  (
  .D(_0334_),
  .CK(clk),
  .Q(\d_pipe[10][14] ),
  .QN(_0021_)
);

DFF_X1 \d_pipe[10][15]$_DFFE_PP_  (
  .D(_0335_),
  .CK(clk),
  .Q(\d_pipe[10][15] ),
  .QN(_0022_)
);

DFF_X1 \d_pipe[10][16]$_DFFE_PP_  (
  .D(_0336_),
  .CK(clk),
  .Q(\d_pipe[10][16] ),
  .QN(_0023_)
);

DFF_X1 \d_pipe[10][17]$_DFFE_PP_  (
  .D(_0337_),
  .CK(clk),
  .Q(\d_pipe[10][17] ),
  .QN(_0024_)
);

DFF_X1 \d_pipe[10][18]$_DFFE_PP_  (
  .D(_0338_),
  .CK(clk),
  .Q(\d_pipe[10][18] ),
  .QN(_0025_)
);

DFF_X1 \d_pipe[10][19]$_DFFE_PP_  (
  .D(_0339_),
  .CK(clk),
  .Q(\d_pipe[10][19] ),
  .QN(_0026_)
);

DFF_X1 \d_pipe[10][20]$_DFFE_PP_  (
  .D(_0340_),
  .CK(clk),
  .Q(\d_pipe[10][20] ),
  .QN(_0027_)
);

DFF_X1 \d_pipe[10][21]$_DFFE_PP_  (
  .D(_0341_),
  .CK(clk),
  .Q(\d_pipe[10][21] ),
  .QN(_0028_)
);

DFF_X1 \d_pipe[10][22]$_DFFE_PP_  (
  .D(_0342_),
  .CK(clk),
  .Q(\d_pipe[10][22] ),
  .QN(_0029_)
);

DFF_X1 \d_pipe[10][23]$_DFFE_PP_  (
  .D(_0343_),
  .CK(clk),
  .Q(\d_pipe[10][23] ),
  .QN(_0030_)
);

DFF_X1 \d_pipe[11][12]$_DFFE_PP_  (
  .D(_0344_),
  .CK(clk),
  .Q(\d_pipe[11][12] ),
  .QN(_4285_)
);

DFF_X1 \d_pipe[11][13]$_DFFE_PP_  (
  .D(_0345_),
  .CK(clk),
  .Q(\d_pipe[11][13] ),
  .QN(_4286_)
);

DFF_X1 \d_pipe[11][14]$_DFFE_PP_  (
  .D(_0346_),
  .CK(clk),
  .Q(\d_pipe[11][14] ),
  .QN(_0011_)
);

DFF_X1 \d_pipe[11][15]$_DFFE_PP_  (
  .D(_0347_),
  .CK(clk),
  .Q(\d_pipe[11][15] ),
  .QN(_0012_)
);

DFF_X1 \d_pipe[11][16]$_DFFE_PP_  (
  .D(_0348_),
  .CK(clk),
  .Q(\d_pipe[11][16] ),
  .QN(_0013_)
);

DFF_X1 \d_pipe[11][17]$_DFFE_PP_  (
  .D(_0349_),
  .CK(clk),
  .Q(\d_pipe[11][17] ),
  .QN(_0014_)
);

DFF_X1 \d_pipe[11][18]$_DFFE_PP_  (
  .D(_0350_),
  .CK(clk),
  .Q(\d_pipe[11][18] ),
  .QN(_0015_)
);

DFF_X1 \d_pipe[11][19]$_DFFE_PP_  (
  .D(_0351_),
  .CK(clk),
  .Q(\d_pipe[11][19] ),
  .QN(_0016_)
);

DFF_X1 \d_pipe[11][20]$_DFFE_PP_  (
  .D(_0352_),
  .CK(clk),
  .Q(\d_pipe[11][20] ),
  .QN(_0017_)
);

DFF_X1 \d_pipe[11][21]$_DFFE_PP_  (
  .D(_0353_),
  .CK(clk),
  .Q(\d_pipe[11][21] ),
  .QN(_0018_)
);

DFF_X1 \d_pipe[11][22]$_DFFE_PP_  (
  .D(_0354_),
  .CK(clk),
  .Q(\d_pipe[11][22] ),
  .QN(_0019_)
);

DFF_X1 \d_pipe[11][23]$_DFFE_PP_  (
  .D(_0355_),
  .CK(clk),
  .Q(\d_pipe[11][23] ),
  .QN(_0020_)
);

DFF_X1 \d_pipe[1][12]$_DFFE_PP_  (
  .D(_0248_),
  .CK(clk),
  .Q(\d_pipe[1][12] ),
  .QN(_4216_)
);

DFF_X1 \d_pipe[1][13]$_DFFE_PP_  (
  .D(_0249_),
  .CK(clk),
  .Q(\d_pipe[1][13] ),
  .QN(_4217_)
);

DFF_X1 \d_pipe[1][14]$_DFFE_PP_  (
  .D(_0250_),
  .CK(clk),
  .Q(\d_pipe[1][14] ),
  .QN(_0001_)
);

DFF_X1 \d_pipe[1][15]$_DFFE_PP_  (
  .D(_0251_),
  .CK(clk),
  .Q(\d_pipe[1][15] ),
  .QN(_0002_)
);

DFF_X1 \d_pipe[1][16]$_DFFE_PP_  (
  .D(_0252_),
  .CK(clk),
  .Q(\d_pipe[1][16] ),
  .QN(_0003_)
);

DFF_X1 \d_pipe[1][17]$_DFFE_PP_  (
  .D(_0253_),
  .CK(clk),
  .Q(\d_pipe[1][17] ),
  .QN(_0004_)
);

DFF_X1 \d_pipe[1][18]$_DFFE_PP_  (
  .D(_0254_),
  .CK(clk),
  .Q(\d_pipe[1][18] ),
  .QN(_0005_)
);

DFF_X1 \d_pipe[1][19]$_DFFE_PP_  (
  .D(_0255_),
  .CK(clk),
  .Q(\d_pipe[1][19] ),
  .QN(_0006_)
);

DFF_X1 \d_pipe[1][20]$_DFFE_PP_  (
  .D(_0256_),
  .CK(clk),
  .Q(\d_pipe[1][20] ),
  .QN(_0007_)
);

DFF_X1 \d_pipe[1][21]$_DFFE_PP_  (
  .D(_0257_),
  .CK(clk),
  .Q(\d_pipe[1][21] ),
  .QN(_0008_)
);

DFF_X1 \d_pipe[1][22]$_DFFE_PP_  (
  .D(_0258_),
  .CK(clk),
  .Q(\d_pipe[1][22] ),
  .QN(_0009_)
);

DFF_X1 \d_pipe[1][23]$_DFFE_PP_  (
  .D(_0259_),
  .CK(clk),
  .Q(\d_pipe[1][23] ),
  .QN(_0010_)
);

DFF_X1 \d_pipe[2][12]$_DFFE_PP_  (
  .D(_0169_),
  .CK(clk),
  .Q(\d_pipe[2][12] ),
  .QN(_4144_)
);

DFF_X1 \d_pipe[2][13]$_DFFE_PP_  (
  .D(_0170_),
  .CK(clk),
  .Q(\d_pipe[2][13] ),
  .QN(_4145_)
);

DFF_X1 \d_pipe[2][14]$_DFFE_PP_  (
  .D(_0171_),
  .CK(clk),
  .Q(\d_pipe[2][14] ),
  .QN(_0091_)
);

DFF_X1 \d_pipe[2][15]$_DFFE_PP_  (
  .D(_0172_),
  .CK(clk),
  .Q(\d_pipe[2][15] ),
  .QN(_0092_)
);

DFF_X1 \d_pipe[2][16]$_DFFE_PP_  (
  .D(_0173_),
  .CK(clk),
  .Q(\d_pipe[2][16] ),
  .QN(_0093_)
);

DFF_X1 \d_pipe[2][17]$_DFFE_PP_  (
  .D(_0174_),
  .CK(clk),
  .Q(\d_pipe[2][17] ),
  .QN(_0094_)
);

DFF_X1 \d_pipe[2][18]$_DFFE_PP_  (
  .D(_0175_),
  .CK(clk),
  .Q(\d_pipe[2][18] ),
  .QN(_0095_)
);

DFF_X1 \d_pipe[2][19]$_DFFE_PP_  (
  .D(_0176_),
  .CK(clk),
  .Q(\d_pipe[2][19] ),
  .QN(_0096_)
);

DFF_X1 \d_pipe[2][20]$_DFFE_PP_  (
  .D(_0177_),
  .CK(clk),
  .Q(\d_pipe[2][20] ),
  .QN(_0097_)
);

DFF_X1 \d_pipe[2][21]$_DFFE_PP_  (
  .D(_0178_),
  .CK(clk),
  .Q(\d_pipe[2][21] ),
  .QN(_0098_)
);

DFF_X1 \d_pipe[2][22]$_DFFE_PP_  (
  .D(_0179_),
  .CK(clk),
  .Q(\d_pipe[2][22] ),
  .QN(_0099_)
);

DFF_X1 \d_pipe[2][23]$_DFFE_PP_  (
  .D(_0180_),
  .CK(clk),
  .Q(\d_pipe[2][23] ),
  .QN(_0100_)
);

DFF_X1 \d_pipe[3][12]$_DFFE_PP_  (
  .D(_0157_),
  .CK(clk),
  .Q(\d_pipe[3][12] ),
  .QN(_4180_)
);

DFF_X1 \d_pipe[3][13]$_DFFE_PP_  (
  .D(_0158_),
  .CK(clk),
  .Q(\d_pipe[3][13] ),
  .QN(_4181_)
);

DFF_X1 \d_pipe[3][14]$_DFFE_PP_  (
  .D(_0159_),
  .CK(clk),
  .Q(\d_pipe[3][14] ),
  .QN(_0101_)
);

DFF_X1 \d_pipe[3][15]$_DFFE_PP_  (
  .D(_0160_),
  .CK(clk),
  .Q(\d_pipe[3][15] ),
  .QN(_0102_)
);

DFF_X1 \d_pipe[3][16]$_DFFE_PP_  (
  .D(_0161_),
  .CK(clk),
  .Q(\d_pipe[3][16] ),
  .QN(_0103_)
);

DFF_X1 \d_pipe[3][17]$_DFFE_PP_  (
  .D(_0162_),
  .CK(clk),
  .Q(\d_pipe[3][17] ),
  .QN(_0104_)
);

DFF_X1 \d_pipe[3][18]$_DFFE_PP_  (
  .D(_0163_),
  .CK(clk),
  .Q(\d_pipe[3][18] ),
  .QN(_0105_)
);

DFF_X1 \d_pipe[3][19]$_DFFE_PP_  (
  .D(_0164_),
  .CK(clk),
  .Q(\d_pipe[3][19] ),
  .QN(_0106_)
);

DFF_X1 \d_pipe[3][20]$_DFFE_PP_  (
  .D(_0165_),
  .CK(clk),
  .Q(\d_pipe[3][20] ),
  .QN(_0107_)
);

DFF_X1 \d_pipe[3][21]$_DFFE_PP_  (
  .D(_0166_),
  .CK(clk),
  .Q(\d_pipe[3][21] ),
  .QN(_0108_)
);

DFF_X1 \d_pipe[3][22]$_DFFE_PP_  (
  .D(_0167_),
  .CK(clk),
  .Q(\d_pipe[3][22] ),
  .QN(_0109_)
);

DFF_X1 \d_pipe[3][23]$_DFFE_PP_  (
  .D(_0168_),
  .CK(clk),
  .Q(\d_pipe[3][23] ),
  .QN(_0110_)
);

DFF_X1 \d_pipe[4][12]$_DFFE_PP_  (
  .D(_0260_),
  .CK(clk),
  .Q(\d_pipe[4][12] ),
  .QN(_4537_)
);

DFF_X1 \d_pipe[4][13]$_DFFE_PP_  (
  .D(_0261_),
  .CK(clk),
  .Q(\d_pipe[4][13] ),
  .QN(_4538_)
);

DFF_X1 \d_pipe[4][14]$_DFFE_PP_  (
  .D(_0262_),
  .CK(clk),
  .Q(\d_pipe[4][14] ),
  .QN(_0081_)
);

DFF_X1 \d_pipe[4][15]$_DFFE_PP_  (
  .D(_0263_),
  .CK(clk),
  .Q(\d_pipe[4][15] ),
  .QN(_0082_)
);

DFF_X1 \d_pipe[4][16]$_DFFE_PP_  (
  .D(_0264_),
  .CK(clk),
  .Q(\d_pipe[4][16] ),
  .QN(_0083_)
);

DFF_X1 \d_pipe[4][17]$_DFFE_PP_  (
  .D(_0265_),
  .CK(clk),
  .Q(\d_pipe[4][17] ),
  .QN(_0084_)
);

DFF_X1 \d_pipe[4][18]$_DFFE_PP_  (
  .D(_0266_),
  .CK(clk),
  .Q(\d_pipe[4][18] ),
  .QN(_0085_)
);

DFF_X1 \d_pipe[4][19]$_DFFE_PP_  (
  .D(_0267_),
  .CK(clk),
  .Q(\d_pipe[4][19] ),
  .QN(_0086_)
);

DFF_X1 \d_pipe[4][20]$_DFFE_PP_  (
  .D(_0268_),
  .CK(clk),
  .Q(\d_pipe[4][20] ),
  .QN(_0087_)
);

DFF_X1 \d_pipe[4][21]$_DFFE_PP_  (
  .D(_0269_),
  .CK(clk),
  .Q(\d_pipe[4][21] ),
  .QN(_0088_)
);

DFF_X1 \d_pipe[4][22]$_DFFE_PP_  (
  .D(_0270_),
  .CK(clk),
  .Q(\d_pipe[4][22] ),
  .QN(_0089_)
);

DFF_X1 \d_pipe[4][23]$_DFFE_PP_  (
  .D(_0271_),
  .CK(clk),
  .Q(\d_pipe[4][23] ),
  .QN(_0090_)
);

DFF_X1 \d_pipe[5][12]$_DFFE_PP_  (
  .D(_0272_),
  .CK(clk),
  .Q(\d_pipe[5][12] ),
  .QN(_4501_)
);

DFF_X1 \d_pipe[5][13]$_DFFE_PP_  (
  .D(_0273_),
  .CK(clk),
  .Q(\d_pipe[5][13] ),
  .QN(_4502_)
);

DFF_X1 \d_pipe[5][14]$_DFFE_PP_  (
  .D(_0274_),
  .CK(clk),
  .Q(\d_pipe[5][14] ),
  .QN(_0071_)
);

DFF_X1 \d_pipe[5][15]$_DFFE_PP_  (
  .D(_0275_),
  .CK(clk),
  .Q(\d_pipe[5][15] ),
  .QN(_0072_)
);

DFF_X1 \d_pipe[5][16]$_DFFE_PP_  (
  .D(_0276_),
  .CK(clk),
  .Q(\d_pipe[5][16] ),
  .QN(_0073_)
);

DFF_X1 \d_pipe[5][17]$_DFFE_PP_  (
  .D(_0277_),
  .CK(clk),
  .Q(\d_pipe[5][17] ),
  .QN(_0074_)
);

DFF_X1 \d_pipe[5][18]$_DFFE_PP_  (
  .D(_0278_),
  .CK(clk),
  .Q(\d_pipe[5][18] ),
  .QN(_0075_)
);

DFF_X1 \d_pipe[5][19]$_DFFE_PP_  (
  .D(_0279_),
  .CK(clk),
  .Q(\d_pipe[5][19] ),
  .QN(_0076_)
);

DFF_X1 \d_pipe[5][20]$_DFFE_PP_  (
  .D(_0280_),
  .CK(clk),
  .Q(\d_pipe[5][20] ),
  .QN(_0077_)
);

DFF_X1 \d_pipe[5][21]$_DFFE_PP_  (
  .D(_0281_),
  .CK(clk),
  .Q(\d_pipe[5][21] ),
  .QN(_0078_)
);

DFF_X1 \d_pipe[5][22]$_DFFE_PP_  (
  .D(_0282_),
  .CK(clk),
  .Q(\d_pipe[5][22] ),
  .QN(_0079_)
);

DFF_X1 \d_pipe[5][23]$_DFFE_PP_  (
  .D(_0283_),
  .CK(clk),
  .Q(\d_pipe[5][23] ),
  .QN(_0080_)
);

DFF_X1 \d_pipe[6][12]$_DFFE_PP_  (
  .D(_0284_),
  .CK(clk),
  .Q(\d_pipe[6][12] ),
  .QN(_4465_)
);

DFF_X1 \d_pipe[6][13]$_DFFE_PP_  (
  .D(_0285_),
  .CK(clk),
  .Q(\d_pipe[6][13] ),
  .QN(_4466_)
);

DFF_X1 \d_pipe[6][14]$_DFFE_PP_  (
  .D(_0286_),
  .CK(clk),
  .Q(\d_pipe[6][14] ),
  .QN(_0061_)
);

DFF_X1 \d_pipe[6][15]$_DFFE_PP_  (
  .D(_0287_),
  .CK(clk),
  .Q(\d_pipe[6][15] ),
  .QN(_0062_)
);

DFF_X1 \d_pipe[6][16]$_DFFE_PP_  (
  .D(_0288_),
  .CK(clk),
  .Q(\d_pipe[6][16] ),
  .QN(_0063_)
);

DFF_X1 \d_pipe[6][17]$_DFFE_PP_  (
  .D(_0289_),
  .CK(clk),
  .Q(\d_pipe[6][17] ),
  .QN(_0064_)
);

DFF_X1 \d_pipe[6][18]$_DFFE_PP_  (
  .D(_0290_),
  .CK(clk),
  .Q(\d_pipe[6][18] ),
  .QN(_0065_)
);

DFF_X1 \d_pipe[6][19]$_DFFE_PP_  (
  .D(_0291_),
  .CK(clk),
  .Q(\d_pipe[6][19] ),
  .QN(_0066_)
);

DFF_X1 \d_pipe[6][20]$_DFFE_PP_  (
  .D(_0292_),
  .CK(clk),
  .Q(\d_pipe[6][20] ),
  .QN(_0067_)
);

DFF_X1 \d_pipe[6][21]$_DFFE_PP_  (
  .D(_0293_),
  .CK(clk),
  .Q(\d_pipe[6][21] ),
  .QN(_0068_)
);

DFF_X1 \d_pipe[6][22]$_DFFE_PP_  (
  .D(_0294_),
  .CK(clk),
  .Q(\d_pipe[6][22] ),
  .QN(_0069_)
);

DFF_X1 \d_pipe[6][23]$_DFFE_PP_  (
  .D(_0295_),
  .CK(clk),
  .Q(\d_pipe[6][23] ),
  .QN(_0070_)
);

DFF_X1 \d_pipe[7][12]$_DFFE_PP_  (
  .D(_0296_),
  .CK(clk),
  .Q(\d_pipe[7][12] ),
  .QN(_4429_)
);

DFF_X1 \d_pipe[7][13]$_DFFE_PP_  (
  .D(_0297_),
  .CK(clk),
  .Q(\d_pipe[7][13] ),
  .QN(_4430_)
);

DFF_X1 \d_pipe[7][14]$_DFFE_PP_  (
  .D(_0298_),
  .CK(clk),
  .Q(\d_pipe[7][14] ),
  .QN(_0051_)
);

DFF_X1 \d_pipe[7][15]$_DFFE_PP_  (
  .D(_0299_),
  .CK(clk),
  .Q(\d_pipe[7][15] ),
  .QN(_0052_)
);

DFF_X1 \d_pipe[7][16]$_DFFE_PP_  (
  .D(_0300_),
  .CK(clk),
  .Q(\d_pipe[7][16] ),
  .QN(_0053_)
);

DFF_X1 \d_pipe[7][17]$_DFFE_PP_  (
  .D(_0301_),
  .CK(clk),
  .Q(\d_pipe[7][17] ),
  .QN(_0054_)
);

DFF_X1 \d_pipe[7][18]$_DFFE_PP_  (
  .D(_0302_),
  .CK(clk),
  .Q(\d_pipe[7][18] ),
  .QN(_0055_)
);

DFF_X1 \d_pipe[7][19]$_DFFE_PP_  (
  .D(_0303_),
  .CK(clk),
  .Q(\d_pipe[7][19] ),
  .QN(_0056_)
);

DFF_X1 \d_pipe[7][20]$_DFFE_PP_  (
  .D(_0304_),
  .CK(clk),
  .Q(\d_pipe[7][20] ),
  .QN(_0057_)
);

DFF_X1 \d_pipe[7][21]$_DFFE_PP_  (
  .D(_0305_),
  .CK(clk),
  .Q(\d_pipe[7][21] ),
  .QN(_0058_)
);

DFF_X1 \d_pipe[7][22]$_DFFE_PP_  (
  .D(_0306_),
  .CK(clk),
  .Q(\d_pipe[7][22] ),
  .QN(_0059_)
);

DFF_X1 \d_pipe[7][23]$_DFFE_PP_  (
  .D(_0307_),
  .CK(clk),
  .Q(\d_pipe[7][23] ),
  .QN(_0060_)
);

DFF_X1 \d_pipe[8][12]$_DFFE_PP_  (
  .D(_0308_),
  .CK(clk),
  .Q(\d_pipe[8][12] ),
  .QN(_4393_)
);

DFF_X1 \d_pipe[8][13]$_DFFE_PP_  (
  .D(_0309_),
  .CK(clk),
  .Q(\d_pipe[8][13] ),
  .QN(_4394_)
);

DFF_X1 \d_pipe[8][14]$_DFFE_PP_  (
  .D(_0310_),
  .CK(clk),
  .Q(\d_pipe[8][14] ),
  .QN(_0041_)
);

DFF_X1 \d_pipe[8][15]$_DFFE_PP_  (
  .D(_0311_),
  .CK(clk),
  .Q(\d_pipe[8][15] ),
  .QN(_0042_)
);

DFF_X1 \d_pipe[8][16]$_DFFE_PP_  (
  .D(_0312_),
  .CK(clk),
  .Q(\d_pipe[8][16] ),
  .QN(_0043_)
);

DFF_X1 \d_pipe[8][17]$_DFFE_PP_  (
  .D(_0313_),
  .CK(clk),
  .Q(\d_pipe[8][17] ),
  .QN(_0044_)
);

DFF_X1 \d_pipe[8][18]$_DFFE_PP_  (
  .D(_0314_),
  .CK(clk),
  .Q(\d_pipe[8][18] ),
  .QN(_0045_)
);

DFF_X1 \d_pipe[8][19]$_DFFE_PP_  (
  .D(_0315_),
  .CK(clk),
  .Q(\d_pipe[8][19] ),
  .QN(_0046_)
);

DFF_X1 \d_pipe[8][20]$_DFFE_PP_  (
  .D(_0316_),
  .CK(clk),
  .Q(\d_pipe[8][20] ),
  .QN(_0047_)
);

DFF_X1 \d_pipe[8][21]$_DFFE_PP_  (
  .D(_0317_),
  .CK(clk),
  .Q(\d_pipe[8][21] ),
  .QN(_0048_)
);

DFF_X1 \d_pipe[8][22]$_DFFE_PP_  (
  .D(_0318_),
  .CK(clk),
  .Q(\d_pipe[8][22] ),
  .QN(_0049_)
);

DFF_X1 \d_pipe[8][23]$_DFFE_PP_  (
  .D(_0319_),
  .CK(clk),
  .Q(\d_pipe[8][23] ),
  .QN(_0050_)
);

DFF_X1 \d_pipe[9][12]$_DFFE_PP_  (
  .D(_0320_),
  .CK(clk),
  .Q(\d_pipe[9][12] ),
  .QN(_4357_)
);

DFF_X1 \q[0]$_DFFE_PP_  (
  .D(_0210_),
  .CK(clk),
  .Q(q[0]),
  .QN(_4002_)
);

DFF_X1 \q[10]$_DFFE_PP_  (
  .D(_0220_),
  .CK(clk),
  .Q(q[10]),
  .QN(_3992_)
);

DFF_X1 \q[11]$_DFFE_PP_  (
  .D(_0221_),
  .CK(clk),
  .Q(q[11]),
  .QN(_3991_)
);

DFF_X1 \q[1]$_DFFE_PP_  (
  .D(_0211_),
  .CK(clk),
  .Q(q[1]),
  .QN(_4001_)
);

DFF_X1 \q[2]$_DFFE_PP_  (
  .D(_0212_),
  .CK(clk),
  .Q(q[2]),
  .QN(_4000_)
);

DFF_X1 \q[3]$_DFFE_PP_  (
  .D(_0213_),
  .CK(clk),
  .Q(q[3]),
  .QN(_3999_)
);

DFF_X1 \q[4]$_DFFE_PP_  (
  .D(_0214_),
  .CK(clk),
  .Q(q[4]),
  .QN(_3998_)
);

DFF_X1 \q[5]$_DFFE_PP_  (
  .D(_0215_),
  .CK(clk),
  .Q(q[5]),
  .QN(_3997_)
);

DFF_X1 \q[6]$_DFFE_PP_  (
  .D(_0216_),
  .CK(clk),
  .Q(q[6]),
  .QN(_3996_)
);

DFF_X1 \q[7]$_DFFE_PP_  (
  .D(_0217_),
  .CK(clk),
  .Q(q[7]),
  .QN(_3995_)
);

DFF_X1 \q[8]$_DFFE_PP_  (
  .D(_0218_),
  .CK(clk),
  .Q(q[8]),
  .QN(_3994_)
);

DFF_X1 \q[9]$_DFFE_PP_  (
  .D(_0219_),
  .CK(clk),
  .Q(q[9]),
  .QN(_3993_)
);

DFF_X1 \q_pipe[10][0]$_DFFE_PP_  (
  .D(_0562_),
  .CK(clk),
  .Q(\q_pipe[10][0] ),
  .QN(_3774_)
);

DFF_X1 \q_pipe[10][1]$_DFFE_PP_  (
  .D(_0563_),
  .CK(clk),
  .Q(\q_pipe[10][1] ),
  .QN(_3773_)
);

DFF_X1 \q_pipe[10][2]$_DFFE_PP_  (
  .D(_0564_),
  .CK(clk),
  .Q(\q_pipe[10][2] ),
  .QN(_3772_)
);

DFF_X1 \q_pipe[10][3]$_DFFE_PP_  (
  .D(_0565_),
  .CK(clk),
  .Q(\q_pipe[10][3] ),
  .QN(_3771_)
);

DFF_X1 \q_pipe[10][4]$_DFFE_PP_  (
  .D(_0566_),
  .CK(clk),
  .Q(\q_pipe[10][4] ),
  .QN(_3770_)
);

DFF_X1 \q_pipe[10][5]$_DFFE_PP_  (
  .D(_0567_),
  .CK(clk),
  .Q(\q_pipe[10][5] ),
  .QN(_3769_)
);

DFF_X1 \q_pipe[10][6]$_DFFE_PP_  (
  .D(_0568_),
  .CK(clk),
  .Q(\q_pipe[10][6] ),
  .QN(_3768_)
);

DFF_X1 \q_pipe[10][7]$_DFFE_PP_  (
  .D(_0569_),
  .CK(clk),
  .Q(\q_pipe[10][7] ),
  .QN(_3767_)
);

DFF_X1 \q_pipe[10][8]$_DFFE_PP_  (
  .D(_0570_),
  .CK(clk),
  .Q(\q_pipe[10][8] ),
  .QN(_3766_)
);

DFF_X1 \q_pipe[10][9]$_DFFE_PP_  (
  .D(_0571_),
  .CK(clk),
  .Q(\q_pipe[10][9] ),
  .QN(_3765_)
);

DFF_X1 \q_pipe[11][0]$_DFFE_PP_  (
  .D(_0572_),
  .CK(clk),
  .Q(\q_pipe[11][0] ),
  .QN(_3764_)
);

DFF_X1 \q_pipe[11][10]$_DFFE_PP_  (
  .D(_0582_),
  .CK(clk),
  .Q(\q_pipe[11][10] ),
  .QN(_3754_)
);

DFF_X1 \q_pipe[11][1]$_DFFE_PP_  (
  .D(_0573_),
  .CK(clk),
  .Q(\q_pipe[11][1] ),
  .QN(_3763_)
);

DFF_X1 \q_pipe[11][2]$_DFFE_PP_  (
  .D(_0574_),
  .CK(clk),
  .Q(\q_pipe[11][2] ),
  .QN(_3762_)
);

DFF_X1 \q_pipe[11][3]$_DFFE_PP_  (
  .D(_0575_),
  .CK(clk),
  .Q(\q_pipe[11][3] ),
  .QN(_3761_)
);

DFF_X1 \q_pipe[11][4]$_DFFE_PP_  (
  .D(_0576_),
  .CK(clk),
  .Q(\q_pipe[11][4] ),
  .QN(_3760_)
);

DFF_X1 \q_pipe[11][5]$_DFFE_PP_  (
  .D(_0577_),
  .CK(clk),
  .Q(\q_pipe[11][5] ),
  .QN(_3759_)
);

DFF_X1 \q_pipe[11][6]$_DFFE_PP_  (
  .D(_0578_),
  .CK(clk),
  .Q(\q_pipe[11][6] ),
  .QN(_3758_)
);

DFF_X1 \q_pipe[11][7]$_DFFE_PP_  (
  .D(_0579_),
  .CK(clk),
  .Q(\q_pipe[11][7] ),
  .QN(_3757_)
);

DFF_X1 \q_pipe[11][8]$_DFFE_PP_  (
  .D(_0580_),
  .CK(clk),
  .Q(\q_pipe[11][8] ),
  .QN(_3756_)
);

DFF_X1 \q_pipe[11][9]$_DFFE_PP_  (
  .D(_0581_),
  .CK(clk),
  .Q(\q_pipe[11][9] ),
  .QN(_3755_)
);

DFF_X1 \q_pipe[1]$_DFFE_PP_  (
  .D(_0209_),
  .CK(clk),
  .Q(\q_pipe[1] ),
  .QN(_4003_)
);

DFF_X1 \q_pipe[2][0]$_DFFE_PP_  (
  .D(_0518_),
  .CK(clk),
  .Q(\q_pipe[2][0] ),
  .QN(_3818_)
);

DFF_X1 \q_pipe[2][1]$_DFFE_PP_  (
  .D(_0519_),
  .CK(clk),
  .Q(\q_pipe[2][1] ),
  .QN(_3817_)
);

DFF_X1 \q_pipe[3][0]$_DFFE_PP_  (
  .D(_0520_),
  .CK(clk),
  .Q(\q_pipe[3][0] ),
  .QN(_3816_)
);

DFF_X1 \q_pipe[3][1]$_DFFE_PP_  (
  .D(_0521_),
  .CK(clk),
  .Q(\q_pipe[3][1] ),
  .QN(_3815_)
);

DFF_X1 \q_pipe[3][2]$_DFFE_PP_  (
  .D(_0522_),
  .CK(clk),
  .Q(\q_pipe[3][2] ),
  .QN(_3814_)
);

DFF_X1 \q_pipe[4][0]$_DFFE_PP_  (
  .D(_0523_),
  .CK(clk),
  .Q(\q_pipe[4][0] ),
  .QN(_3813_)
);

DFF_X1 \q_pipe[4][1]$_DFFE_PP_  (
  .D(_0524_),
  .CK(clk),
  .Q(\q_pipe[4][1] ),
  .QN(_3812_)
);

DFF_X1 \q_pipe[4][2]$_DFFE_PP_  (
  .D(_0525_),
  .CK(clk),
  .Q(\q_pipe[4][2] ),
  .QN(_3811_)
);

DFF_X1 \q_pipe[4][3]$_DFFE_PP_  (
  .D(_0526_),
  .CK(clk),
  .Q(\q_pipe[4][3] ),
  .QN(_3810_)
);

DFF_X1 \q_pipe[5][0]$_DFFE_PP_  (
  .D(_0527_),
  .CK(clk),
  .Q(\q_pipe[5][0] ),
  .QN(_3809_)
);

DFF_X1 \q_pipe[5][1]$_DFFE_PP_  (
  .D(_0528_),
  .CK(clk),
  .Q(\q_pipe[5][1] ),
  .QN(_3808_)
);

DFF_X1 \q_pipe[5][2]$_DFFE_PP_  (
  .D(_0529_),
  .CK(clk),
  .Q(\q_pipe[5][2] ),
  .QN(_3807_)
);

DFF_X1 \q_pipe[5][3]$_DFFE_PP_  (
  .D(_0530_),
  .CK(clk),
  .Q(\q_pipe[5][3] ),
  .QN(_3806_)
);

DFF_X1 \q_pipe[5][4]$_DFFE_PP_  (
  .D(_0531_),
  .CK(clk),
  .Q(\q_pipe[5][4] ),
  .QN(_3805_)
);

DFF_X1 \q_pipe[6][0]$_DFFE_PP_  (
  .D(_0532_),
  .CK(clk),
  .Q(\q_pipe[6][0] ),
  .QN(_3804_)
);

DFF_X1 \q_pipe[6][1]$_DFFE_PP_  (
  .D(_0533_),
  .CK(clk),
  .Q(\q_pipe[6][1] ),
  .QN(_3803_)
);

DFF_X1 \q_pipe[6][2]$_DFFE_PP_  (
  .D(_0534_),
  .CK(clk),
  .Q(\q_pipe[6][2] ),
  .QN(_3802_)
);

DFF_X1 \q_pipe[6][3]$_DFFE_PP_  (
  .D(_0535_),
  .CK(clk),
  .Q(\q_pipe[6][3] ),
  .QN(_3801_)
);

DFF_X1 \q_pipe[6][4]$_DFFE_PP_  (
  .D(_0536_),
  .CK(clk),
  .Q(\q_pipe[6][4] ),
  .QN(_3800_)
);

DFF_X1 \q_pipe[6][5]$_DFFE_PP_  (
  .D(_0537_),
  .CK(clk),
  .Q(\q_pipe[6][5] ),
  .QN(_3799_)
);

DFF_X1 \q_pipe[7][0]$_DFFE_PP_  (
  .D(_0538_),
  .CK(clk),
  .Q(\q_pipe[7][0] ),
  .QN(_3798_)
);

DFF_X1 \q_pipe[7][1]$_DFFE_PP_  (
  .D(_0539_),
  .CK(clk),
  .Q(\q_pipe[7][1] ),
  .QN(_3797_)
);

DFF_X1 \q_pipe[7][2]$_DFFE_PP_  (
  .D(_0540_),
  .CK(clk),
  .Q(\q_pipe[7][2] ),
  .QN(_3796_)
);

DFF_X1 \q_pipe[7][3]$_DFFE_PP_  (
  .D(_0541_),
  .CK(clk),
  .Q(\q_pipe[7][3] ),
  .QN(_3795_)
);

DFF_X1 \q_pipe[7][4]$_DFFE_PP_  (
  .D(_0542_),
  .CK(clk),
  .Q(\q_pipe[7][4] ),
  .QN(_3794_)
);

DFF_X1 \q_pipe[7][5]$_DFFE_PP_  (
  .D(_0543_),
  .CK(clk),
  .Q(\q_pipe[7][5] ),
  .QN(_3793_)
);

DFF_X1 \q_pipe[7][6]$_DFFE_PP_  (
  .D(_0544_),
  .CK(clk),
  .Q(\q_pipe[7][6] ),
  .QN(_3792_)
);

DFF_X1 \q_pipe[8][0]$_DFFE_PP_  (
  .D(_0545_),
  .CK(clk),
  .Q(\q_pipe[8][0] ),
  .QN(_3791_)
);

DFF_X1 \q_pipe[8][1]$_DFFE_PP_  (
  .D(_0546_),
  .CK(clk),
  .Q(\q_pipe[8][1] ),
  .QN(_3790_)
);

DFF_X1 \q_pipe[8][2]$_DFFE_PP_  (
  .D(_0547_),
  .CK(clk),
  .Q(\q_pipe[8][2] ),
  .QN(_3789_)
);

DFF_X1 \q_pipe[8][3]$_DFFE_PP_  (
  .D(_0548_),
  .CK(clk),
  .Q(\q_pipe[8][3] ),
  .QN(_3788_)
);

DFF_X1 \q_pipe[8][4]$_DFFE_PP_  (
  .D(_0549_),
  .CK(clk),
  .Q(\q_pipe[8][4] ),
  .QN(_3787_)
);

DFF_X1 \q_pipe[8][5]$_DFFE_PP_  (
  .D(_0550_),
  .CK(clk),
  .Q(\q_pipe[8][5] ),
  .QN(_3786_)
);

DFF_X1 \q_pipe[8][6]$_DFFE_PP_  (
  .D(_0551_),
  .CK(clk),
  .Q(\q_pipe[8][6] ),
  .QN(_3785_)
);

DFF_X1 \q_pipe[8][7]$_DFFE_PP_  (
  .D(_0552_),
  .CK(clk),
  .Q(\q_pipe[8][7] ),
  .QN(_3784_)
);

DFF_X1 \q_pipe[9]$_DFFE_PP_  (
  .D(_0553_),
  .CK(clk),
  .Q(\q_pipe[9] ),
  .QN(_3783_)
);

DFF_X1 \s_pipe[10][10]$_DFFE_PP_  (
  .D(_0503_),
  .CK(clk),
  .Q(\s_pipe[10][10] ),
  .QN(_3831_)
);

DFF_X1 \s_pipe[10][11]$_DFFE_PP_  (
  .D(_0504_),
  .CK(clk),
  .Q(\s_pipe[10][11] ),
  .QN(_3830_)
);

DFF_X1 \s_pipe[10][12]$_DFFE_PP_  (
  .D(_0505_),
  .CK(clk),
  .Q(\s_pipe[10][12] ),
  .QN(_4073_)
);

DFF_X1 \s_pipe[10][13]$_DFFE_PP_  (
  .D(_0506_),
  .CK(clk),
  .Q(\s_pipe[10][13] ),
  .QN(_3829_)
);

DFF_X1 \s_pipe[10][14]$_DFFE_PP_  (
  .D(_0507_),
  .CK(clk),
  .Q(\s_pipe[10][14] ),
  .QN(_3828_)
);

DFF_X1 \s_pipe[10][15]$_DFFE_PP_  (
  .D(_0508_),
  .CK(clk),
  .Q(\s_pipe[10][15] ),
  .QN(_3827_)
);

DFF_X1 \s_pipe[10][16]$_DFFE_PP_  (
  .D(_0509_),
  .CK(clk),
  .Q(\s_pipe[10][16] ),
  .QN(_3826_)
);

DFF_X1 \s_pipe[10][17]$_DFFE_PP_  (
  .D(_0510_),
  .CK(clk),
  .Q(\s_pipe[10][17] ),
  .QN(_3825_)
);

DFF_X1 \s_pipe[10][18]$_DFFE_PP_  (
  .D(_0511_),
  .CK(clk),
  .Q(\s_pipe[10][18] ),
  .QN(_3824_)
);

DFF_X1 \s_pipe[10][19]$_DFFE_PP_  (
  .D(_0512_),
  .CK(clk),
  .Q(\s_pipe[10][19] ),
  .QN(_3823_)
);

DFF_X1 \s_pipe[10][20]$_DFFE_PP_  (
  .D(_0513_),
  .CK(clk),
  .Q(\s_pipe[10][20] ),
  .QN(_3822_)
);

DFF_X1 \s_pipe[10][21]$_DFFE_PP_  (
  .D(_0514_),
  .CK(clk),
  .Q(\s_pipe[10][21] ),
  .QN(_3821_)
);

DFF_X1 \s_pipe[10][22]$_DFFE_PP_  (
  .D(_0515_),
  .CK(clk),
  .Q(\s_pipe[10][22] ),
  .QN(_3820_)
);

DFF_X1 \s_pipe[10][23]$_DFFE_PP_  (
  .D(_0516_),
  .CK(clk),
  .Q(\s_pipe[10][23] ),
  .QN(_3819_)
);

DFF_X1 \s_pipe[10][24]$_DFFE_PP_  (
  .D(_0517_),
  .CK(clk),
  .Q(\s_pipe[10][24] ),
  .QN(_0120_)
);

DFF_X1 \s_pipe[11][11]$_DFFE_PP_  (
  .D(_0413_),
  .CK(clk),
  .Q(\s_pipe[11][11] ),
  .QN(_3911_)
);

DFF_X1 \s_pipe[11][12]$_DFFE_PP_  (
  .D(_0414_),
  .CK(clk),
  .Q(\s_pipe[11][12] ),
  .QN(_4066_)
);

DFF_X1 \s_pipe[11][13]$_DFFE_PP_  (
  .D(_0415_),
  .CK(clk),
  .Q(\s_pipe[11][13] ),
  .QN(_3910_)
);

DFF_X1 \s_pipe[11][14]$_DFFE_PP_  (
  .D(_0416_),
  .CK(clk),
  .Q(\s_pipe[11][14] ),
  .QN(_3909_)
);

DFF_X1 \s_pipe[11][15]$_DFFE_PP_  (
  .D(_0417_),
  .CK(clk),
  .Q(\s_pipe[11][15] ),
  .QN(_3908_)
);

DFF_X1 \s_pipe[11][16]$_DFFE_PP_  (
  .D(_0418_),
  .CK(clk),
  .Q(\s_pipe[11][16] ),
  .QN(_3907_)
);

DFF_X1 \s_pipe[11][17]$_DFFE_PP_  (
  .D(_0419_),
  .CK(clk),
  .Q(\s_pipe[11][17] ),
  .QN(_3906_)
);

DFF_X1 \s_pipe[11][18]$_DFFE_PP_  (
  .D(_0420_),
  .CK(clk),
  .Q(\s_pipe[11][18] ),
  .QN(_3905_)
);

DFF_X1 \s_pipe[11][19]$_DFFE_PP_  (
  .D(_0421_),
  .CK(clk),
  .Q(\s_pipe[11][19] ),
  .QN(_3904_)
);

DFF_X1 \s_pipe[11][20]$_DFFE_PP_  (
  .D(_0422_),
  .CK(clk),
  .Q(\s_pipe[11][20] ),
  .QN(_3903_)
);

DFF_X1 \s_pipe[11][21]$_DFFE_PP_  (
  .D(_0423_),
  .CK(clk),
  .Q(\s_pipe[11][21] ),
  .QN(_3902_)
);

DFF_X1 \s_pipe[11][22]$_DFFE_PP_  (
  .D(_0424_),
  .CK(clk),
  .Q(\s_pipe[11][22] ),
  .QN(_3901_)
);

DFF_X1 \s_pipe[11][23]$_DFFE_PP_  (
  .D(_0425_),
  .CK(clk),
  .Q(\s_pipe[11][23] ),
  .QN(_3900_)
);

DFF_X1 \s_pipe[11][24]$_DFFE_PP_  (
  .D(_0426_),
  .CK(clk),
  .Q(\s_pipe[11][24] ),
  .QN(_0121_)
);

DFF_X1 \s_pipe[12][24]$_DFFE_PP_  (
  .D(_0156_),
  .CK(clk),
  .Q(\s_pipe[12][24] ),
  .QN(_0122_)
);

DFF_X1 \s_pipe[1][10]$_DFFE_PP_  (
  .D(_0190_),
  .CK(clk),
  .Q(\s_pipe[1][10] ),
  .QN(_4020_)
);

DFF_X1 \s_pipe[1][11]$_DFFE_PP_  (
  .D(_0191_),
  .CK(clk),
  .Q(\s_pipe[1][11] ),
  .QN(_4019_)
);

DFF_X1 \s_pipe[1][12]$_DFFE_PP_  (
  .D(_0192_),
  .CK(clk),
  .Q(\s_pipe[1][12] ),
  .QN(_4056_)
);

DFF_X1 \s_pipe[1][13]$_DFFE_PP_  (
  .D(_0193_),
  .CK(clk),
  .Q(\s_pipe[1][13] ),
  .QN(_4018_)
);

DFF_X1 \s_pipe[1][14]$_DFFE_PP_  (
  .D(_0194_),
  .CK(clk),
  .Q(\s_pipe[1][14] ),
  .QN(_4017_)
);

DFF_X1 \s_pipe[1][15]$_DFFE_PP_  (
  .D(_0195_),
  .CK(clk),
  .Q(\s_pipe[1][15] ),
  .QN(_4016_)
);

DFF_X1 \s_pipe[1][16]$_DFFE_PP_  (
  .D(_0196_),
  .CK(clk),
  .Q(\s_pipe[1][16] ),
  .QN(_4015_)
);

DFF_X1 \s_pipe[1][17]$_DFFE_PP_  (
  .D(_0197_),
  .CK(clk),
  .Q(\s_pipe[1][17] ),
  .QN(_4014_)
);

DFF_X1 \s_pipe[1][18]$_DFFE_PP_  (
  .D(_0198_),
  .CK(clk),
  .Q(\s_pipe[1][18] ),
  .QN(_4013_)
);

DFF_X1 \s_pipe[1][19]$_DFFE_PP_  (
  .D(_0199_),
  .CK(clk),
  .Q(\s_pipe[1][19] ),
  .QN(_4012_)
);

DFF_X1 \s_pipe[1][1]$_DFFE_PP_  (
  .D(_0181_),
  .CK(clk),
  .Q(\s_pipe[1][1] ),
  .QN(_4029_)
);

DFF_X1 \s_pipe[1][20]$_DFFE_PP_  (
  .D(_0200_),
  .CK(clk),
  .Q(\s_pipe[1][20] ),
  .QN(_4011_)
);

DFF_X1 \s_pipe[1][21]$_DFFE_PP_  (
  .D(_0201_),
  .CK(clk),
  .Q(\s_pipe[1][21] ),
  .QN(_4010_)
);

DFF_X1 \s_pipe[1][22]$_DFFE_PP_  (
  .D(_0202_),
  .CK(clk),
  .Q(\s_pipe[1][22] ),
  .QN(_4009_)
);

DFF_X1 \s_pipe[1][23]$_DFFE_PP_  (
  .D(_0203_),
  .CK(clk),
  .Q(\s_pipe[1][23] ),
  .QN(_4008_)
);

DFF_X1 \s_pipe[1][24]$_DFFE_PP_  (
  .D(_0204_),
  .CK(clk),
  .Q(\s_pipe[1][24] ),
  .QN(_0111_)
);

DFF_X1 \s_pipe[1][2]$_DFFE_PP_  (
  .D(_0182_),
  .CK(clk),
  .Q(\s_pipe[1][2] ),
  .QN(_4028_)
);

DFF_X1 \s_pipe[1][3]$_DFFE_PP_  (
  .D(_0183_),
  .CK(clk),
  .Q(\s_pipe[1][3] ),
  .QN(_4027_)
);

DFF_X1 \s_pipe[1][4]$_DFFE_PP_  (
  .D(_0184_),
  .CK(clk),
  .Q(\s_pipe[1][4] ),
  .QN(_4026_)
);

DFF_X1 \s_pipe[1][5]$_DFFE_PP_  (
  .D(_0185_),
  .CK(clk),
  .Q(\s_pipe[1][5] ),
  .QN(_4025_)
);

DFF_X1 \s_pipe[1][6]$_DFFE_PP_  (
  .D(_0186_),
  .CK(clk),
  .Q(\s_pipe[1][6] ),
  .QN(_4024_)
);

DFF_X1 \s_pipe[1][7]$_DFFE_PP_  (
  .D(_0187_),
  .CK(clk),
  .Q(\s_pipe[1][7] ),
  .QN(_4023_)
);

DFF_X1 \s_pipe[1][8]$_DFFE_PP_  (
  .D(_0188_),
  .CK(clk),
  .Q(\s_pipe[1][8] ),
  .QN(_4022_)
);

DFF_X1 \s_pipe[1][9]$_DFFE_PP_  (
  .D(_0189_),
  .CK(clk),
  .Q(\s_pipe[1][9] ),
  .QN(_4021_)
);

DFF_X1 \s_pipe[2][10]$_DFFE_PP_  (
  .D(_0376_),
  .CK(clk),
  .Q(\s_pipe[2][10] ),
  .QN(_3944_)
);

DFF_X1 \s_pipe[2][11]$_DFFE_PP_  (
  .D(_0377_),
  .CK(clk),
  .Q(\s_pipe[2][11] ),
  .QN(_3943_)
);

DFF_X1 \s_pipe[2][12]$_DFFE_PP_  (
  .D(_0378_),
  .CK(clk),
  .Q(\s_pipe[2][12] ),
  .QN(_4042_)
);

DFF_X1 \s_pipe[2][13]$_DFFE_PP_  (
  .D(_0379_),
  .CK(clk),
  .Q(\s_pipe[2][13] ),
  .QN(_3942_)
);

DFF_X1 \s_pipe[2][14]$_DFFE_PP_  (
  .D(_0380_),
  .CK(clk),
  .Q(\s_pipe[2][14] ),
  .QN(_3941_)
);

DFF_X1 \s_pipe[2][15]$_DFFE_PP_  (
  .D(_0381_),
  .CK(clk),
  .Q(\s_pipe[2][15] ),
  .QN(_3940_)
);

DFF_X1 \s_pipe[2][16]$_DFFE_PP_  (
  .D(_0382_),
  .CK(clk),
  .Q(\s_pipe[2][16] ),
  .QN(_3939_)
);

DFF_X1 \s_pipe[2][17]$_DFFE_PP_  (
  .D(_0383_),
  .CK(clk),
  .Q(\s_pipe[2][17] ),
  .QN(_3938_)
);

DFF_X1 \s_pipe[2][18]$_DFFE_PP_  (
  .D(_0384_),
  .CK(clk),
  .Q(\s_pipe[2][18] ),
  .QN(_3937_)
);

DFF_X1 \s_pipe[2][19]$_DFFE_PP_  (
  .D(_0385_),
  .CK(clk),
  .Q(\s_pipe[2][19] ),
  .QN(_3936_)
);

DFF_X1 \s_pipe[2][20]$_DFFE_PP_  (
  .D(_0386_),
  .CK(clk),
  .Q(\s_pipe[2][20] ),
  .QN(_3935_)
);

DFF_X1 \s_pipe[2][21]$_DFFE_PP_  (
  .D(_0387_),
  .CK(clk),
  .Q(\s_pipe[2][21] ),
  .QN(_3934_)
);

DFF_X1 \s_pipe[2][22]$_DFFE_PP_  (
  .D(_0388_),
  .CK(clk),
  .Q(\s_pipe[2][22] ),
  .QN(_3933_)
);

DFF_X1 \s_pipe[2][23]$_DFFE_PP_  (
  .D(_0389_),
  .CK(clk),
  .Q(\s_pipe[2][23] ),
  .QN(_3932_)
);

DFF_X1 \s_pipe[2][24]$_DFFE_PP_  (
  .D(_0390_),
  .CK(clk),
  .Q(\s_pipe[2][24] ),
  .QN(_0112_)
);

DFF_X1 \s_pipe[2][2]$_DFFE_PP_  (
  .D(_0368_),
  .CK(clk),
  .Q(\s_pipe[2][2] ),
  .QN(_3952_)
);

DFF_X1 \s_pipe[2][3]$_DFFE_PP_  (
  .D(_0369_),
  .CK(clk),
  .Q(\s_pipe[2][3] ),
  .QN(_3951_)
);

DFF_X1 \s_pipe[2][4]$_DFFE_PP_  (
  .D(_0370_),
  .CK(clk),
  .Q(\s_pipe[2][4] ),
  .QN(_3950_)
);

DFF_X1 \s_pipe[2][5]$_DFFE_PP_  (
  .D(_0371_),
  .CK(clk),
  .Q(\s_pipe[2][5] ),
  .QN(_3949_)
);

DFF_X1 \s_pipe[2][6]$_DFFE_PP_  (
  .D(_0372_),
  .CK(clk),
  .Q(\s_pipe[2][6] ),
  .QN(_3948_)
);

DFF_X1 \s_pipe[2][7]$_DFFE_PP_  (
  .D(_0373_),
  .CK(clk),
  .Q(\s_pipe[2][7] ),
  .QN(_3947_)
);

DFF_X1 \s_pipe[2][8]$_DFFE_PP_  (
  .D(_0374_),
  .CK(clk),
  .Q(\s_pipe[2][8] ),
  .QN(_3946_)
);

DFF_X1 \s_pipe[2][9]$_DFFE_PP_  (
  .D(_0375_),
  .CK(clk),
  .Q(\s_pipe[2][9] ),
  .QN(_3945_)
);

DFF_X1 \s_pipe[3][10]$_DFFE_PP_  (
  .D(_0398_),
  .CK(clk),
  .Q(\s_pipe[3][10] ),
  .QN(_3924_)
);

DFF_X1 \s_pipe[3][11]$_DFFE_PP_  (
  .D(_0399_),
  .CK(clk),
  .Q(\s_pipe[3][11] ),
  .QN(_3923_)
);

DFF_X1 \s_pipe[3][12]$_DFFE_PP_  (
  .D(_0400_),
  .CK(clk),
  .Q(\s_pipe[3][12] ),
  .QN(_4049_)
);

DFF_X1 \s_pipe[3][13]$_DFFE_PP_  (
  .D(_0401_),
  .CK(clk),
  .Q(\s_pipe[3][13] ),
  .QN(_3922_)
);

DFF_X1 \s_pipe[3][14]$_DFFE_PP_  (
  .D(_0402_),
  .CK(clk),
  .Q(\s_pipe[3][14] ),
  .QN(_3921_)
);

DFF_X1 \s_pipe[3][15]$_DFFE_PP_  (
  .D(_0403_),
  .CK(clk),
  .Q(\s_pipe[3][15] ),
  .QN(_3920_)
);

DFF_X1 \s_pipe[3][16]$_DFFE_PP_  (
  .D(_0404_),
  .CK(clk),
  .Q(\s_pipe[3][16] ),
  .QN(_3919_)
);

DFF_X1 \s_pipe[3][17]$_DFFE_PP_  (
  .D(_0405_),
  .CK(clk),
  .Q(\s_pipe[3][17] ),
  .QN(_3918_)
);

DFF_X1 \s_pipe[3][18]$_DFFE_PP_  (
  .D(_0406_),
  .CK(clk),
  .Q(\s_pipe[3][18] ),
  .QN(_3917_)
);

DFF_X1 \s_pipe[3][19]$_DFFE_PP_  (
  .D(_0407_),
  .CK(clk),
  .Q(\s_pipe[3][19] ),
  .QN(_3916_)
);

DFF_X1 \s_pipe[3][20]$_DFFE_PP_  (
  .D(_0408_),
  .CK(clk),
  .Q(\s_pipe[3][20] ),
  .QN(_3915_)
);

DFF_X1 \s_pipe[3][21]$_DFFE_PP_  (
  .D(_0409_),
  .CK(clk),
  .Q(\s_pipe[3][21] ),
  .QN(_3914_)
);

DFF_X1 \s_pipe[3][22]$_DFFE_PP_  (
  .D(_0410_),
  .CK(clk),
  .Q(\s_pipe[3][22] ),
  .QN(_3913_)
);

DFF_X1 \s_pipe[3][23]$_DFFE_PP_  (
  .D(_0411_),
  .CK(clk),
  .Q(\s_pipe[3][23] ),
  .QN(_3912_)
);

DFF_X1 \s_pipe[3][24]$_DFFE_PP_  (
  .D(_0412_),
  .CK(clk),
  .Q(\s_pipe[3][24] ),
  .QN(_0113_)
);

DFF_X1 \s_pipe[3][3]$_DFFE_PP_  (
  .D(_0391_),
  .CK(clk),
  .Q(\s_pipe[3][3] ),
  .QN(_3931_)
);

DFF_X1 \s_pipe[3][4]$_DFFE_PP_  (
  .D(_0392_),
  .CK(clk),
  .Q(\s_pipe[3][4] ),
  .QN(_3930_)
);

DFF_X1 \s_pipe[3][5]$_DFFE_PP_  (
  .D(_0393_),
  .CK(clk),
  .Q(\s_pipe[3][5] ),
  .QN(_3929_)
);

DFF_X1 \s_pipe[3][6]$_DFFE_PP_  (
  .D(_0394_),
  .CK(clk),
  .Q(\s_pipe[3][6] ),
  .QN(_3928_)
);

DFF_X1 \s_pipe[3][7]$_DFFE_PP_  (
  .D(_0395_),
  .CK(clk),
  .Q(\s_pipe[3][7] ),
  .QN(_3927_)
);

DFF_X1 \s_pipe[3][8]$_DFFE_PP_  (
  .D(_0396_),
  .CK(clk),
  .Q(\s_pipe[3][8] ),
  .QN(_3926_)
);

DFF_X1 \s_pipe[3][9]$_DFFE_PP_  (
  .D(_0397_),
  .CK(clk),
  .Q(\s_pipe[3][9] ),
  .QN(_3925_)
);

DFF_X1 \s_pipe[4][10]$_DFFE_PP_  (
  .D(_0433_),
  .CK(clk),
  .Q(\s_pipe[4][10] ),
  .QN(_3893_)
);

DFF_X1 \s_pipe[4][11]$_DFFE_PP_  (
  .D(_0434_),
  .CK(clk),
  .Q(\s_pipe[4][11] ),
  .QN(_3892_)
);

DFF_X1 \s_pipe[4][12]$_DFFE_PP_  (
  .D(_0435_),
  .CK(clk),
  .Q(\s_pipe[4][12] ),
  .QN(_4115_)
);

DFF_X1 \s_pipe[4][13]$_DFFE_PP_  (
  .D(_0436_),
  .CK(clk),
  .Q(\s_pipe[4][13] ),
  .QN(_3891_)
);

DFF_X1 \s_pipe[4][14]$_DFFE_PP_  (
  .D(_0437_),
  .CK(clk),
  .Q(\s_pipe[4][14] ),
  .QN(_3890_)
);

DFF_X1 \s_pipe[4][15]$_DFFE_PP_  (
  .D(_0438_),
  .CK(clk),
  .Q(\s_pipe[4][15] ),
  .QN(_3889_)
);

DFF_X1 \s_pipe[4][16]$_DFFE_PP_  (
  .D(_0439_),
  .CK(clk),
  .Q(\s_pipe[4][16] ),
  .QN(_3888_)
);

DFF_X1 \s_pipe[4][17]$_DFFE_PP_  (
  .D(_0440_),
  .CK(clk),
  .Q(\s_pipe[4][17] ),
  .QN(_3887_)
);

DFF_X1 \s_pipe[4][18]$_DFFE_PP_  (
  .D(_0441_),
  .CK(clk),
  .Q(\s_pipe[4][18] ),
  .QN(_3886_)
);

DFF_X1 \s_pipe[4][19]$_DFFE_PP_  (
  .D(_0442_),
  .CK(clk),
  .Q(\s_pipe[4][19] ),
  .QN(_3885_)
);

DFF_X1 \s_pipe[4][20]$_DFFE_PP_  (
  .D(_0443_),
  .CK(clk),
  .Q(\s_pipe[4][20] ),
  .QN(_3884_)
);

DFF_X1 \s_pipe[4][21]$_DFFE_PP_  (
  .D(_0444_),
  .CK(clk),
  .Q(\s_pipe[4][21] ),
  .QN(_3883_)
);

DFF_X1 \s_pipe[4][22]$_DFFE_PP_  (
  .D(_0445_),
  .CK(clk),
  .Q(\s_pipe[4][22] ),
  .QN(_3882_)
);

DFF_X1 \s_pipe[4][23]$_DFFE_PP_  (
  .D(_0446_),
  .CK(clk),
  .Q(\s_pipe[4][23] ),
  .QN(_3881_)
);

DFF_X1 \s_pipe[4][24]$_DFFE_PP_  (
  .D(_0447_),
  .CK(clk),
  .Q(\s_pipe[4][24] ),
  .QN(_0114_)
);

DFF_X1 \s_pipe[4][4]$_DFFE_PP_  (
  .D(_0427_),
  .CK(clk),
  .Q(\s_pipe[4][4] ),
  .QN(_3899_)
);

DFF_X1 \s_pipe[4][5]$_DFFE_PP_  (
  .D(_0428_),
  .CK(clk),
  .Q(\s_pipe[4][5] ),
  .QN(_3898_)
);

DFF_X1 \s_pipe[4][6]$_DFFE_PP_  (
  .D(_0429_),
  .CK(clk),
  .Q(\s_pipe[4][6] ),
  .QN(_3897_)
);

DFF_X1 \s_pipe[4][7]$_DFFE_PP_  (
  .D(_0430_),
  .CK(clk),
  .Q(\s_pipe[4][7] ),
  .QN(_3896_)
);

DFF_X1 \s_pipe[4][8]$_DFFE_PP_  (
  .D(_0431_),
  .CK(clk),
  .Q(\s_pipe[4][8] ),
  .QN(_3895_)
);

DFF_X1 \s_pipe[4][9]$_DFFE_PP_  (
  .D(_0432_),
  .CK(clk),
  .Q(\s_pipe[4][9] ),
  .QN(_3894_)
);

DFF_X1 \s_pipe[5][10]$_DFFE_PP_  (
  .D(_0469_),
  .CK(clk),
  .Q(\s_pipe[5][10] ),
  .QN(_3861_)
);

DFF_X1 \s_pipe[5][11]$_DFFE_PP_  (
  .D(_0470_),
  .CK(clk),
  .Q(\s_pipe[5][11] ),
  .QN(_3860_)
);

DFF_X1 \s_pipe[5][12]$_DFFE_PP_  (
  .D(_0471_),
  .CK(clk),
  .Q(\s_pipe[5][12] ),
  .QN(_4108_)
);

DFF_X1 \s_pipe[5][13]$_DFFE_PP_  (
  .D(_0472_),
  .CK(clk),
  .Q(\s_pipe[5][13] ),
  .QN(_3859_)
);

DFF_X1 \s_pipe[5][14]$_DFFE_PP_  (
  .D(_0473_),
  .CK(clk),
  .Q(\s_pipe[5][14] ),
  .QN(_3858_)
);

DFF_X1 \s_pipe[5][15]$_DFFE_PP_  (
  .D(_0474_),
  .CK(clk),
  .Q(\s_pipe[5][15] ),
  .QN(_3857_)
);

DFF_X1 \s_pipe[5][16]$_DFFE_PP_  (
  .D(_0475_),
  .CK(clk),
  .Q(\s_pipe[5][16] ),
  .QN(_3856_)
);

DFF_X1 \s_pipe[5][17]$_DFFE_PP_  (
  .D(_0476_),
  .CK(clk),
  .Q(\s_pipe[5][17] ),
  .QN(_3855_)
);

DFF_X1 \s_pipe[5][18]$_DFFE_PP_  (
  .D(_0477_),
  .CK(clk),
  .Q(\s_pipe[5][18] ),
  .QN(_3854_)
);

DFF_X1 \s_pipe[5][19]$_DFFE_PP_  (
  .D(_0478_),
  .CK(clk),
  .Q(\s_pipe[5][19] ),
  .QN(_3853_)
);

DFF_X1 \s_pipe[5][20]$_DFFE_PP_  (
  .D(_0479_),
  .CK(clk),
  .Q(\s_pipe[5][20] ),
  .QN(_3852_)
);

DFF_X1 \s_pipe[5][21]$_DFFE_PP_  (
  .D(_0480_),
  .CK(clk),
  .Q(\s_pipe[5][21] ),
  .QN(_3851_)
);

DFF_X1 \s_pipe[5][22]$_DFFE_PP_  (
  .D(_0481_),
  .CK(clk),
  .Q(\s_pipe[5][22] ),
  .QN(_3850_)
);

DFF_X1 \s_pipe[5][23]$_DFFE_PP_  (
  .D(_0482_),
  .CK(clk),
  .Q(\s_pipe[5][23] ),
  .QN(_3849_)
);

DFF_X1 \s_pipe[5][24]$_DFFE_PP_  (
  .D(_0483_),
  .CK(clk),
  .Q(\s_pipe[5][24] ),
  .QN(_0115_)
);

DFF_X1 \s_pipe[5][5]$_DFFE_PP_  (
  .D(_0464_),
  .CK(clk),
  .Q(\s_pipe[5][5] ),
  .QN(_3866_)
);

DFF_X1 \s_pipe[5][6]$_DFFE_PP_  (
  .D(_0465_),
  .CK(clk),
  .Q(\s_pipe[5][6] ),
  .QN(_3865_)
);

DFF_X1 \s_pipe[5][7]$_DFFE_PP_  (
  .D(_0466_),
  .CK(clk),
  .Q(\s_pipe[5][7] ),
  .QN(_3864_)
);

DFF_X1 \s_pipe[5][8]$_DFFE_PP_  (
  .D(_0467_),
  .CK(clk),
  .Q(\s_pipe[5][8] ),
  .QN(_3863_)
);

DFF_X1 \s_pipe[5][9]$_DFFE_PP_  (
  .D(_0468_),
  .CK(clk),
  .Q(\s_pipe[5][9] ),
  .QN(_3862_)
);

DFF_X1 \s_pipe[6][10]$_DFFE_PP_  (
  .D(_0488_),
  .CK(clk),
  .Q(\s_pipe[6][10] ),
  .QN(_3844_)
);

DFF_X1 \s_pipe[6][11]$_DFFE_PP_  (
  .D(_0489_),
  .CK(clk),
  .Q(\s_pipe[6][11] ),
  .QN(_3843_)
);

DFF_X1 \s_pipe[6][12]$_DFFE_PP_  (
  .D(_0490_),
  .CK(clk),
  .Q(\s_pipe[6][12] ),
  .QN(_4101_)
);

DFF_X1 \s_pipe[6][13]$_DFFE_PP_  (
  .D(_0491_),
  .CK(clk),
  .Q(\s_pipe[6][13] ),
  .QN(_3842_)
);

DFF_X1 \s_pipe[6][14]$_DFFE_PP_  (
  .D(_0492_),
  .CK(clk),
  .Q(\s_pipe[6][14] ),
  .QN(_3841_)
);

DFF_X1 \s_pipe[6][15]$_DFFE_PP_  (
  .D(_0493_),
  .CK(clk),
  .Q(\s_pipe[6][15] ),
  .QN(_3840_)
);

DFF_X1 \s_pipe[6][16]$_DFFE_PP_  (
  .D(_0494_),
  .CK(clk),
  .Q(\s_pipe[6][16] ),
  .QN(_3839_)
);

DFF_X1 \s_pipe[6][17]$_DFFE_PP_  (
  .D(_0495_),
  .CK(clk),
  .Q(\s_pipe[6][17] ),
  .QN(_3838_)
);

DFF_X1 \s_pipe[6][18]$_DFFE_PP_  (
  .D(_0496_),
  .CK(clk),
  .Q(\s_pipe[6][18] ),
  .QN(_3837_)
);

DFF_X1 \s_pipe[6][19]$_DFFE_PP_  (
  .D(_0497_),
  .CK(clk),
  .Q(\s_pipe[6][19] ),
  .QN(_3836_)
);

DFF_X1 \s_pipe[6][20]$_DFFE_PP_  (
  .D(_0498_),
  .CK(clk),
  .Q(\s_pipe[6][20] ),
  .QN(_3835_)
);

DFF_X1 \s_pipe[6][21]$_DFFE_PP_  (
  .D(_0499_),
  .CK(clk),
  .Q(\s_pipe[6][21] ),
  .QN(_3834_)
);

DFF_X1 \s_pipe[6][22]$_DFFE_PP_  (
  .D(_0500_),
  .CK(clk),
  .Q(\s_pipe[6][22] ),
  .QN(_3833_)
);

DFF_X1 \s_pipe[6][23]$_DFFE_PP_  (
  .D(_0501_),
  .CK(clk),
  .Q(\s_pipe[6][23] ),
  .QN(_3832_)
);

DFF_X1 \s_pipe[6][24]$_DFFE_PP_  (
  .D(_0502_),
  .CK(clk),
  .Q(\s_pipe[6][24] ),
  .QN(_0116_)
);

DFF_X1 \s_pipe[6][6]$_DFFE_PP_  (
  .D(_0484_),
  .CK(clk),
  .Q(\s_pipe[6][6] ),
  .QN(_3848_)
);

DFF_X1 \s_pipe[6][7]$_DFFE_PP_  (
  .D(_0485_),
  .CK(clk),
  .Q(\s_pipe[6][7] ),
  .QN(_3847_)
);

DFF_X1 \s_pipe[6][8]$_DFFE_PP_  (
  .D(_0486_),
  .CK(clk),
  .Q(\s_pipe[6][8] ),
  .QN(_3846_)
);

DFF_X1 \s_pipe[6][9]$_DFFE_PP_  (
  .D(_0487_),
  .CK(clk),
  .Q(\s_pipe[6][9] ),
  .QN(_3845_)
);

DFF_X1 \s_pipe[7][10]$_DFFE_PP_  (
  .D(_0586_),
  .CK(clk),
  .Q(\s_pipe[7][10] ),
  .QN(_3750_)
);

DFF_X1 \s_pipe[7][11]$_DFFE_PP_  (
  .D(_0587_),
  .CK(clk),
  .Q(\s_pipe[7][11] ),
  .QN(_3749_)
);

DFF_X1 \s_pipe[7][12]$_DFFE_PP_  (
  .D(_0588_),
  .CK(clk),
  .Q(\s_pipe[7][12] ),
  .QN(_4094_)
);

DFF_X1 \s_pipe[7][13]$_DFFE_PP_  (
  .D(_0589_),
  .CK(clk),
  .Q(\s_pipe[7][13] ),
  .QN(_3748_)
);

DFF_X1 \s_pipe[7][14]$_DFFE_PP_  (
  .D(_0590_),
  .CK(clk),
  .Q(\s_pipe[7][14] ),
  .QN(_3747_)
);

DFF_X1 \s_pipe[7][15]$_DFFE_PP_  (
  .D(_0591_),
  .CK(clk),
  .Q(\s_pipe[7][15] ),
  .QN(_3746_)
);

DFF_X1 \s_pipe[7][16]$_DFFE_PP_  (
  .D(_0592_),
  .CK(clk),
  .Q(\s_pipe[7][16] ),
  .QN(_3745_)
);

DFF_X1 \s_pipe[7][17]$_DFFE_PP_  (
  .D(_0593_),
  .CK(clk),
  .Q(\s_pipe[7][17] ),
  .QN(_3744_)
);

DFF_X1 \s_pipe[7][18]$_DFFE_PP_  (
  .D(_0594_),
  .CK(clk),
  .Q(\s_pipe[7][18] ),
  .QN(_3743_)
);

DFF_X1 \s_pipe[7][19]$_DFFE_PP_  (
  .D(_0595_),
  .CK(clk),
  .Q(\s_pipe[7][19] ),
  .QN(_3742_)
);

DFF_X1 \s_pipe[7][20]$_DFFE_PP_  (
  .D(_0596_),
  .CK(clk),
  .Q(\s_pipe[7][20] ),
  .QN(_3741_)
);

DFF_X1 \s_pipe[7][21]$_DFFE_PP_  (
  .D(_0597_),
  .CK(clk),
  .Q(\s_pipe[7][21] ),
  .QN(_3740_)
);

DFF_X1 \s_pipe[7][22]$_DFFE_PP_  (
  .D(_0598_),
  .CK(clk),
  .Q(\s_pipe[7][22] ),
  .QN(_3739_)
);

DFF_X1 \s_pipe[7][23]$_DFFE_PP_  (
  .D(_0599_),
  .CK(clk),
  .Q(\s_pipe[7][23] ),
  .QN(_3738_)
);

DFF_X1 \s_pipe[7][24]$_DFFE_PP_  (
  .D(_0600_),
  .CK(clk),
  .Q(\s_pipe[7][24] ),
  .QN(_0117_)
);

DFF_X1 \s_pipe[7][7]$_DFFE_PP_  (
  .D(_0583_),
  .CK(clk),
  .Q(\s_pipe[7][7] ),
  .QN(_3753_)
);

DFF_X1 \s_pipe[7][8]$_DFFE_PP_  (
  .D(_0584_),
  .CK(clk),
  .Q(\s_pipe[7][8] ),
  .QN(_3752_)
);

DFF_X1 \s_pipe[7][9]$_DFFE_PP_  (
  .D(_0585_),
  .CK(clk),
  .Q(\s_pipe[7][9] ),
  .QN(_3751_)
);

DFF_X1 \s_pipe[8][10]$_DFFE_PP_  (
  .D(_0603_),
  .CK(clk),
  .Q(\s_pipe[8][10] ),
  .QN(_3735_)
);

DFF_X1 \s_pipe[8][11]$_DFFE_PP_  (
  .D(_0604_),
  .CK(clk),
  .Q(\s_pipe[8][11] ),
  .QN(_3734_)
);

DFF_X1 \s_pipe[8][12]$_DFFE_PP_  (
  .D(_0605_),
  .CK(clk),
  .Q(\s_pipe[8][12] ),
  .QN(_4087_)
);

DFF_X1 \s_pipe[8][13]$_DFFE_PP_  (
  .D(_0606_),
  .CK(clk),
  .Q(\s_pipe[8][13] ),
  .QN(_3733_)
);

DFF_X1 \s_pipe[8][14]$_DFFE_PP_  (
  .D(_0607_),
  .CK(clk),
  .Q(\s_pipe[8][14] ),
  .QN(_3732_)
);

DFF_X1 \s_pipe[8][15]$_DFFE_PP_  (
  .D(_0608_),
  .CK(clk),
  .Q(\s_pipe[8][15] ),
  .QN(_3731_)
);

DFF_X1 \s_pipe[8][16]$_DFFE_PP_  (
  .D(_0609_),
  .CK(clk),
  .Q(\s_pipe[8][16] ),
  .QN(_3730_)
);

DFF_X1 \s_pipe[8][17]$_DFFE_PP_  (
  .D(_0610_),
  .CK(clk),
  .Q(\s_pipe[8][17] ),
  .QN(_3729_)
);

DFF_X1 \s_pipe[8][18]$_DFFE_PP_  (
  .D(_0611_),
  .CK(clk),
  .Q(\s_pipe[8][18] ),
  .QN(_3728_)
);

DFF_X1 \s_pipe[8][19]$_DFFE_PP_  (
  .D(_0612_),
  .CK(clk),
  .Q(\s_pipe[8][19] ),
  .QN(_3727_)
);

DFF_X1 \s_pipe[8][20]$_DFFE_PP_  (
  .D(_0613_),
  .CK(clk),
  .Q(\s_pipe[8][20] ),
  .QN(_3726_)
);

DFF_X1 \s_pipe[8][21]$_DFFE_PP_  (
  .D(_0614_),
  .CK(clk),
  .Q(\s_pipe[8][21] ),
  .QN(_3725_)
);

DFF_X1 \s_pipe[8][22]$_DFFE_PP_  (
  .D(_0615_),
  .CK(clk),
  .Q(\s_pipe[8][22] ),
  .QN(_3724_)
);

DFF_X1 \s_pipe[8][23]$_DFFE_PP_  (
  .D(_0616_),
  .CK(clk),
  .Q(\s_pipe[8][23] ),
  .QN(_3723_)
);

DFF_X1 \s_pipe[8][24]$_DFFE_PP_  (
  .D(_0617_),
  .CK(clk),
  .Q(\s_pipe[8][24] ),
  .QN(_0118_)
);

DFF_X1 \s_pipe[8][8]$_DFFE_PP_  (
  .D(_0601_),
  .CK(clk),
  .Q(\s_pipe[8][8] ),
  .QN(_3737_)
);

DFF_X1 \s_pipe[8][9]$_DFFE_PP_  (
  .D(_0602_),
  .CK(clk),
  .Q(\s_pipe[8][9] ),
  .QN(_3736_)
);

DFF_X1 \s_pipe[9][10]$_DFFE_PP_  (
  .D(_0449_),
  .CK(clk),
  .Q(\s_pipe[9][10] ),
  .QN(_3879_)
);

DFF_X1 \s_pipe[9][11]$_DFFE_PP_  (
  .D(_0450_),
  .CK(clk),
  .Q(\s_pipe[9][11] ),
  .QN(_3878_)
);

DFF_X1 \s_pipe[9][12]$_DFFE_PP_  (
  .D(_0451_),
  .CK(clk),
  .Q(\s_pipe[9][12] ),
  .QN(_4080_)
);

DFF_X1 \s_pipe[9][13]$_DFFE_PP_  (
  .D(_0452_),
  .CK(clk),
  .Q(\s_pipe[9][13] ),
  .QN(_3877_)
);

DFF_X1 \s_pipe[9][14]$_DFFE_PP_  (
  .D(_0453_),
  .CK(clk),
  .Q(\s_pipe[9][14] ),
  .QN(_3876_)
);

DFF_X1 \s_pipe[9][9]$_DFFE_PP_  (
  .D(_0448_),
  .CK(clk),
  .Q(\s_pipe[9][9] ),
  .QN(_3880_)
);
endmodule //$paramod$ee2aa8736952ca7eee7f4751cab786a479da4583\div_uu

module \$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac (input clk, input ena,
 input dclr, input [7:0] din, input [10:0] coef, output [21:0] result);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire _0032_;
wire _0033_;
wire _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire _0066_;
wire _0067_;
wire _0068_;
wire _0069_;
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
wire _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
wire _0444_;
wire _0445_;
wire _0446_;
wire _0447_;
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire _0658_;
wire _0659_;
wire _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire _0673_;
wire _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire _0679_;
wire _0680_;
wire _0681_;
wire _0682_;
wire _0683_;
wire _0684_;
wire _0685_;
wire _0686_;
wire _0687_;
wire _0688_;
wire _0689_;
wire _0690_;
wire _0691_;
wire _0692_;
wire _0693_;
wire _0694_;
wire _0695_;
wire _0696_;
wire _0697_;
wire _0698_;
wire _0699_;
wire _0700_;
wire _0701_;
wire _0702_;
wire _0703_;
wire _0704_;
wire _0705_;
wire _0706_;
wire _0707_;
wire _0708_;
wire _0709_;
wire _0710_;
wire _0711_;
wire _0712_;
wire _0713_;
wire _0714_;
wire _0715_;
wire _0716_;
wire _0717_;
wire _0718_;
wire _0719_;
wire _0720_;
wire _0721_;
wire _0722_;
wire _0723_;
wire _0724_;
wire _0725_;
wire _0726_;
wire _0727_;
wire _0728_;
wire _0729_;
wire _0730_;
wire _0731_;
wire _0732_;
wire _0733_;
wire _0734_;
wire _0735_;
wire _0736_;
wire _0737_;
wire _0738_;
wire _0739_;
wire _0740_;
wire _0741_;
wire _0742_;
wire _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0748_;
wire _0749_;
wire _0750_;
wire _0751_;
wire _0752_;
wire _0753_;
wire _0754_;
wire _0755_;
wire _0756_;
wire _0757_;
wire _0758_;
wire _0759_;
wire _0760_;
wire _0761_;
wire _0762_;
wire _0763_;
wire _0764_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire _0780_;
wire _0781_;
wire _0782_;
wire _0783_;
wire _0784_;
wire _0785_;
wire _0786_;
wire _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire _0795_;
wire _0796_;
wire _0797_;
wire _0798_;
wire _0799_;
wire _0800_;
wire _0801_;
wire _0802_;
wire _0803_;
wire _0804_;
wire _0805_;
wire _0806_;
wire _0807_;
wire _0808_;
wire _0809_;
wire _0810_;
wire _0811_;
wire _0812_;
wire _0813_;
wire _0814_;
wire _0815_;
wire _0816_;
wire _0817_;
wire _0818_;
wire _0819_;
wire _0820_;
wire _0821_;
wire _0822_;
wire _0823_;
wire _0824_;
wire _0825_;
wire _0826_;
wire _0827_;
wire _0828_;
wire _0829_;
wire _0830_;
wire _0831_;
wire _0832_;
wire _0833_;
wire _0834_;
wire _0835_;
wire _0836_;
wire _0837_;
wire _0838_;
wire _0839_;
wire _0840_;
wire _0841_;
wire _0842_;
wire _0843_;
wire _0844_;
wire _0845_;
wire _0846_;
wire _0847_;
wire _0848_;
wire _0849_;
wire _0850_;
wire _0851_;
wire _0852_;
wire _0853_;
wire _0854_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0858_;
wire _0859_;
wire _0860_;
wire _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0865_;
wire _0866_;
wire _0867_;
wire _0868_;
wire _0869_;
wire _0870_;
wire _0871_;
wire _0872_;
wire _0873_;
wire _0874_;
wire _0875_;
wire _0876_;
wire _0877_;
wire _0878_;
wire _0879_;
wire _0880_;
wire _0881_;
wire _0882_;
wire _0883_;
wire _0884_;
wire _0885_;
wire _0886_;
wire _0887_;
wire _0888_;
wire _0889_;
wire _0890_;
wire _0891_;
wire _0892_;
wire _0893_;
wire _0894_;
wire _0895_;
wire _0896_;
wire _0897_;
wire _0898_;
wire _0899_;
wire _0900_;
wire _0901_;
wire _0902_;
wire _0903_;
wire _0904_;
wire _0905_;
wire _0906_;
wire _0907_;
wire _0908_;
wire _0909_;
wire _0910_;
wire _0911_;
wire _0912_;
wire _0913_;
wire _0914_;
wire _0915_;
wire _0916_;
wire _0917_;
wire _0918_;
wire _0919_;
wire _0920_;
wire _0921_;
wire _0922_;
wire _0923_;
wire _0924_;
wire _0925_;
wire _0926_;
wire _0927_;
wire _0928_;
wire _0929_;
wire _0930_;
wire _0931_;
wire _0932_;
wire _0933_;
wire _0934_;
wire _0935_;
wire _0936_;
wire _0937_;
wire _0938_;
wire _0939_;
wire _0940_;
wire _0941_;
wire _0942_;
wire _0943_;
wire _0944_;
wire _0945_;
wire _0946_;
wire _0947_;
wire _0948_;
wire _0949_;
wire _0950_;
wire _0951_;
wire _0952_;
wire _0953_;
wire _0954_;
wire _0955_;
wire _0956_;
wire _0957_;
wire _0958_;
wire _0959_;
wire _0960_;
wire _0961_;
wire _0962_;
wire _0963_;
wire _0964_;
wire _0965_;
wire _0966_;
wire _0967_;
wire _0968_;
wire _0969_;
wire _0970_;
wire _0971_;
wire _0972_;
wire _0973_;
wire _0974_;
wire _0975_;
wire _0976_;
wire _0977_;
wire _0978_;
wire _0979_;
wire _0980_;
wire _0981_;
wire _0982_;
wire _0983_;
wire _0984_;
wire _0985_;
wire _0986_;
wire _0987_;
wire _0988_;
wire _0989_;
wire _0990_;
wire _0991_;
wire _0992_;
wire _0993_;
wire _0994_;
wire _0995_;
wire _0996_;
wire _0997_;
wire _0998_;
wire _0999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire \ext_mult_res[0] ;
wire \ext_mult_res[10] ;
wire \ext_mult_res[11] ;
wire \ext_mult_res[12] ;
wire \ext_mult_res[13] ;
wire \ext_mult_res[14] ;
wire \ext_mult_res[15] ;
wire \ext_mult_res[16] ;
wire \ext_mult_res[17] ;
wire \ext_mult_res[18] ;
wire \ext_mult_res[1] ;
wire \ext_mult_res[2] ;
wire \ext_mult_res[3] ;
wire \ext_mult_res[4] ;
wire \ext_mult_res[5] ;
wire \ext_mult_res[6] ;
wire \ext_mult_res[7] ;
wire \ext_mult_res[8] ;
wire \ext_mult_res[9] ;

BUF_X1 _1235_ (
  .A(din[0]),
  .Z(_0326_)
);

BUF_X1 _1236_ (
  .A(coef[1]),
  .Z(_0327_)
);

NAND2_X1 _1237_ (
  .A1(_0326_),
  .A2(_0327_),
  .ZN(_0328_)
);

INV_X1 _1238_ (
  .A(_0328_),
  .ZN(_1130_)
);

CLKBUF_X3 _1239_ (
  .A(coef[0]),
  .Z(_0329_)
);

NAND2_X1 _1240_ (
  .A1(_0329_),
  .A2(din[1]),
  .ZN(_0330_)
);

INV_X1 _1241_ (
  .A(_0330_),
  .ZN(_1131_)
);

BUF_X1 _1242_ (
  .A(coef[2]),
  .Z(_0331_)
);

NAND2_X1 _1243_ (
  .A1(_0326_),
  .A2(_0331_),
  .ZN(_0332_)
);

INV_X1 _1244_ (
  .A(_0332_),
  .ZN(_0681_)
);

BUF_X1 _1245_ (
  .A(din[1]),
  .Z(_0333_)
);

NAND2_X1 _1246_ (
  .A1(_0327_),
  .A2(_0333_),
  .ZN(_0334_)
);

INV_X1 _1247_ (
  .A(_0334_),
  .ZN(_0682_)
);

NAND2_X1 _1248_ (
  .A1(_0329_),
  .A2(din[2]),
  .ZN(_0335_)
);

INV_X1 _1249_ (
  .A(_0335_),
  .ZN(_0683_)
);

BUF_X1 _1250_ (
  .A(coef[3]),
  .Z(_0336_)
);

NAND2_X1 _1251_ (
  .A1(_0326_),
  .A2(_0336_),
  .ZN(_0337_)
);

INV_X1 _1252_ (
  .A(_0337_),
  .ZN(_0686_)
);

NAND2_X1 _1253_ (
  .A1(_0333_),
  .A2(_0331_),
  .ZN(_0338_)
);

INV_X1 _1254_ (
  .A(_0338_),
  .ZN(_0687_)
);

BUF_X1 _1255_ (
  .A(din[2]),
  .Z(_0339_)
);

NAND2_X1 _1256_ (
  .A1(_0327_),
  .A2(_0339_),
  .ZN(_0340_)
);

INV_X1 _1257_ (
  .A(_0340_),
  .ZN(_0688_)
);

BUF_X1 _1258_ (
  .A(din[3]),
  .Z(_0341_)
);

NAND2_X1 _1259_ (
  .A1(_0329_),
  .A2(_0341_),
  .ZN(_0342_)
);

INV_X1 _1260_ (
  .A(_0342_),
  .ZN(_0691_)
);

BUF_X1 _1261_ (
  .A(coef[4]),
  .Z(_0343_)
);

NAND2_X1 _1262_ (
  .A1(_0326_),
  .A2(_0343_),
  .ZN(_0694_)
);

NAND2_X1 _1263_ (
  .A1(_0333_),
  .A2(_0336_),
  .ZN(_0695_)
);

NAND2_X1 _1264_ (
  .A1(_0331_),
  .A2(_0339_),
  .ZN(_0696_)
);

NAND2_X1 _1265_ (
  .A1(_0327_),
  .A2(_0341_),
  .ZN(_0344_)
);

INV_X1 _1266_ (
  .A(_0344_),
  .ZN(_1138_)
);

NAND2_X1 _1267_ (
  .A1(_0329_),
  .A2(din[4]),
  .ZN(_0345_)
);

INV_X1 _1268_ (
  .A(_0345_),
  .ZN(_1139_)
);

BUF_X1 _1269_ (
  .A(coef[5]),
  .Z(_0346_)
);

NAND2_X1 _1270_ (
  .A1(_0326_),
  .A2(_0346_),
  .ZN(_0703_)
);

NAND2_X1 _1271_ (
  .A1(_0333_),
  .A2(_0343_),
  .ZN(_0704_)
);

NAND2_X1 _1272_ (
  .A1(_0339_),
  .A2(_0336_),
  .ZN(_0705_)
);

NAND2_X1 _1273_ (
  .A1(_0331_),
  .A2(_0341_),
  .ZN(_0708_)
);

BUF_X1 _1274_ (
  .A(coef[6]),
  .Z(_0347_)
);

NAND2_X1 _1275_ (
  .A1(_0326_),
  .A2(_0347_),
  .ZN(_0720_)
);

NAND2_X1 _1276_ (
  .A1(_0333_),
  .A2(_0346_),
  .ZN(_0721_)
);

NAND2_X1 _1277_ (
  .A1(_0339_),
  .A2(_0343_),
  .ZN(_0722_)
);

NAND2_X1 _1278_ (
  .A1(_0336_),
  .A2(_0341_),
  .ZN(_0725_)
);

BUF_X1 _1279_ (
  .A(din[6]),
  .Z(_0348_)
);

NAND2_X1 _1280_ (
  .A1(_0329_),
  .A2(_0348_),
  .ZN(_0349_)
);

INV_X1 _1281_ (
  .A(_0349_),
  .ZN(_1151_)
);

BUF_X4 _1282_ (
  .A(coef[8]),
  .Z(_0350_)
);

NAND2_X1 _1283_ (
  .A1(_0326_),
  .A2(_0350_),
  .ZN(_0735_)
);

BUF_X4 _1284_ (
  .A(coef[7]),
  .Z(_0351_)
);

NAND2_X1 _1285_ (
  .A1(_0333_),
  .A2(_0351_),
  .ZN(_0736_)
);

NAND2_X1 _1286_ (
  .A1(_0339_),
  .A2(_0347_),
  .ZN(_0737_)
);

NAND2_X1 _1287_ (
  .A1(_0333_),
  .A2(_0347_),
  .ZN(_0352_)
);

INV_X1 _1288_ (
  .A(_0352_),
  .ZN(_0749_)
);

NAND2_X1 _1289_ (
  .A1(_0339_),
  .A2(_0346_),
  .ZN(_0353_)
);

INV_X1 _1290_ (
  .A(_0353_),
  .ZN(_0750_)
);

NAND2_X1 _1291_ (
  .A1(_0341_),
  .A2(_0346_),
  .ZN(_0740_)
);

BUF_X1 _1292_ (
  .A(din[4]),
  .Z(_0354_)
);

NAND2_X1 _1293_ (
  .A1(_0343_),
  .A2(_0354_),
  .ZN(_0741_)
);

BUF_X1 _1294_ (
  .A(din[5]),
  .Z(_0355_)
);

NAND2_X1 _1295_ (
  .A1(_0336_),
  .A2(_0355_),
  .ZN(_0742_)
);

NAND2_X1 _1296_ (
  .A1(_0341_),
  .A2(_0343_),
  .ZN(_0755_)
);

NAND2_X1 _1297_ (
  .A1(_0336_),
  .A2(_0354_),
  .ZN(_0754_)
);

NAND2_X1 _1298_ (
  .A1(_0331_),
  .A2(_0348_),
  .ZN(_0758_)
);

BUF_X8 _1299_ (
  .A(din[7]),
  .Z(_0356_)
);

NAND2_X1 _1300_ (
  .A1(_0327_),
  .A2(_0356_),
  .ZN(_0759_)
);

INV_X1 _1301_ (
  .A(_0759_),
  .ZN(_0763_)
);

NAND2_X4 _1302_ (
  .A1(_0329_),
  .A2(_0356_),
  .ZN(_0760_)
);

INV_X4 _1303_ (
  .A(_0760_),
  .ZN(_0764_)
);

NAND2_X1 _1304_ (
  .A1(_0327_),
  .A2(_0348_),
  .ZN(_0357_)
);

INV_X1 _1305_ (
  .A(_0357_),
  .ZN(_1161_)
);

BUF_X4 _1306_ (
  .A(coef[9]),
  .Z(_0358_)
);

NAND2_X1 _1307_ (
  .A1(_0326_),
  .A2(_0358_),
  .ZN(_0795_)
);

NAND2_X1 _1308_ (
  .A1(_0333_),
  .A2(_0350_),
  .ZN(_0796_)
);

NAND2_X1 _1309_ (
  .A1(_0339_),
  .A2(_0351_),
  .ZN(_0797_)
);

NAND2_X1 _1310_ (
  .A1(_0341_),
  .A2(_0347_),
  .ZN(_0800_)
);

NAND2_X1 _1311_ (
  .A1(_0354_),
  .A2(_0346_),
  .ZN(_0801_)
);

NAND2_X1 _1312_ (
  .A1(_0343_),
  .A2(_0355_),
  .ZN(_0802_)
);

NAND2_X1 _1313_ (
  .A1(_0336_),
  .A2(_0348_),
  .ZN(_0807_)
);

NAND2_X1 _1314_ (
  .A1(_0331_),
  .A2(_0356_),
  .ZN(_0808_)
);

INV_X1 _1315_ (
  .A(_0808_),
  .ZN(_0873_)
);

BUF_X4 _1316_ (
  .A(coef[10]),
  .Z(_0359_)
);

NAND2_X1 _1317_ (
  .A1(_0326_),
  .A2(_0359_),
  .ZN(_0821_)
);

INV_X1 _1318_ (
  .A(_0821_),
  .ZN(_0854_)
);

NAND2_X1 _1319_ (
  .A1(_0339_),
  .A2(_0350_),
  .ZN(_0823_)
);

NAND2_X1 _1320_ (
  .A1(_0341_),
  .A2(_0351_),
  .ZN(_0826_)
);

NAND2_X1 _1321_ (
  .A1(_0354_),
  .A2(_0347_),
  .ZN(_0827_)
);

NAND2_X1 _1322_ (
  .A1(_0346_),
  .A2(_0355_),
  .ZN(_0828_)
);

NAND2_X1 _1323_ (
  .A1(_0343_),
  .A2(_0348_),
  .ZN(_0834_)
);

NAND2_X1 _1324_ (
  .A1(_0333_),
  .A2(_0359_),
  .ZN(_0360_)
);

INV_X1 _1325_ (
  .A(_0360_),
  .ZN(_0852_)
);

NAND2_X1 _1326_ (
  .A1(_0339_),
  .A2(_0358_),
  .ZN(_0361_)
);

INV_X1 _1327_ (
  .A(_0361_),
  .ZN(_0853_)
);

NAND2_X1 _1328_ (
  .A1(_0341_),
  .A2(_0350_),
  .ZN(_0857_)
);

NAND2_X1 _1329_ (
  .A1(_0354_),
  .A2(_0351_),
  .ZN(_0858_)
);

NAND2_X1 _1330_ (
  .A1(_0355_),
  .A2(_0347_),
  .ZN(_0859_)
);

NAND2_X1 _1331_ (
  .A1(_0346_),
  .A2(_0348_),
  .ZN(_0865_)
);

NAND2_X1 _1332_ (
  .A1(_0343_),
  .A2(_0356_),
  .ZN(_0866_)
);

INV_X1 _1333_ (
  .A(_0866_),
  .ZN(_1002_)
);

NAND2_X1 _1334_ (
  .A1(_0339_),
  .A2(_0359_),
  .ZN(_0362_)
);

INV_X1 _1335_ (
  .A(_0362_),
  .ZN(_0882_)
);

NAND2_X1 _1336_ (
  .A1(_0341_),
  .A2(_0358_),
  .ZN(_0885_)
);

NAND2_X1 _1337_ (
  .A1(_0354_),
  .A2(_0350_),
  .ZN(_0886_)
);

NAND2_X1 _1338_ (
  .A1(_0355_),
  .A2(_0351_),
  .ZN(_0887_)
);

NAND2_X1 _1339_ (
  .A1(_0347_),
  .A2(_0348_),
  .ZN(_0894_)
);

NAND2_X1 _1340_ (
  .A1(_0346_),
  .A2(_0356_),
  .ZN(_0895_)
);

INV_X1 _1341_ (
  .A(_0895_),
  .ZN(_1003_)
);

INV_X1 _1342_ (
  .A(_1177_),
  .ZN(_0792_)
);

NAND2_X1 _1343_ (
  .A1(din[3]),
  .A2(_0359_),
  .ZN(_0919_)
);

INV_X1 _1344_ (
  .A(_0919_),
  .ZN(_0951_)
);

NAND2_X1 _1345_ (
  .A1(_0355_),
  .A2(_0350_),
  .ZN(_0921_)
);

NAND2_X1 _1346_ (
  .A1(_0348_),
  .A2(_0351_),
  .ZN(_0927_)
);

NAND2_X1 _1347_ (
  .A1(_0347_),
  .A2(_0356_),
  .ZN(_0928_)
);

INV_X1 _1348_ (
  .A(_0928_),
  .ZN(_1001_)
);

NAND2_X1 _1349_ (
  .A1(_0354_),
  .A2(_0359_),
  .ZN(_0363_)
);

INV_X1 _1350_ (
  .A(_0363_),
  .ZN(_0952_)
);

NAND2_X1 _1351_ (
  .A1(din[5]),
  .A2(_0358_),
  .ZN(_0364_)
);

INV_X1 _1352_ (
  .A(_0364_),
  .ZN(_0953_)
);

NAND2_X1 _1353_ (
  .A1(_0348_),
  .A2(_0350_),
  .ZN(_0959_)
);

NAND2_X2 _1354_ (
  .A1(_0351_),
  .A2(din[7]),
  .ZN(_0960_)
);

INV_X1 _1355_ (
  .A(_0960_),
  .ZN(_1033_)
);

NAND2_X1 _1356_ (
  .A1(_0355_),
  .A2(_0359_),
  .ZN(_0365_)
);

INV_X1 _1357_ (
  .A(_0365_),
  .ZN(_0986_)
);

NAND2_X1 _1358_ (
  .A1(_0348_),
  .A2(_0358_),
  .ZN(_0992_)
);

NAND2_X2 _1359_ (
  .A1(_0350_),
  .A2(din[7]),
  .ZN(_0993_)
);

INV_X1 _1360_ (
  .A(_0993_),
  .ZN(_1022_)
);

NAND2_X2 _1361_ (
  .A1(din[6]),
  .A2(_0359_),
  .ZN(_1052_)
);

INV_X2 _1362_ (
  .A(_1052_),
  .ZN(_1023_)
);

NAND2_X2 _1363_ (
  .A1(_0356_),
  .A2(_0358_),
  .ZN(_1053_)
);

INV_X4 _1364_ (
  .A(_1053_),
  .ZN(_1024_)
);

INV_X1 _1365_ (
  .A(_0987_),
  .ZN(_1027_)
);

INV_X1 _1366_ (
  .A(_0874_),
  .ZN(_0905_)
);

NAND2_X1 _1367_ (
  .A1(_0331_),
  .A2(_0355_),
  .ZN(_0753_)
);

INV_X1 _1368_ (
  .A(_0785_),
  .ZN(_0786_)
);

NAND2_X1 _1369_ (
  .A1(_0336_),
  .A2(_0356_),
  .ZN(_0833_)
);

INV_X1 _1370_ (
  .A(_0875_),
  .ZN(_0969_)
);

NAND2_X1 _1371_ (
  .A1(_0327_),
  .A2(_0354_),
  .ZN(_0709_)
);

NAND2_X1 _1372_ (
  .A1(_0331_),
  .A2(_0354_),
  .ZN(_0726_)
);

NAND2_X1 _1373_ (
  .A1(_0333_),
  .A2(_0358_),
  .ZN(_0822_)
);

INV_X1 _1374_ (
  .A(_0903_),
  .ZN(_0904_)
);

NAND2_X1 _1375_ (
  .A1(_0354_),
  .A2(_0358_),
  .ZN(_0920_)
);

INV_X1 _1376_ (
  .A(_0936_),
  .ZN(_0938_)
);

INV_X1 _1377_ (
  .A(_0968_),
  .ZN(_0970_)
);

INV_X1 _1378_ (
  .A(_1088_),
  .ZN(_0678_)
);

NAND2_X1 _1379_ (
  .A1(_0329_),
  .A2(_0355_),
  .ZN(_0710_)
);

NAND2_X1 _1380_ (
  .A1(_0327_),
  .A2(_0355_),
  .ZN(_0727_)
);

INV_X1 _1381_ (
  .A(_1152_),
  .ZN(_0787_)
);

INV_X1 _1382_ (
  .A(_1186_),
  .ZN(_0879_)
);

INV_X1 _1383_ (
  .A(_1193_),
  .ZN(_0916_)
);

NAND2_X1 _1384_ (
  .A1(_0356_),
  .A2(_0359_),
  .ZN(_1054_)
);

INV_X1 _1385_ (
  .A(_1029_),
  .ZN(_1067_)
);

INV_X1 _1386_ (
  .A(_0752_),
  .ZN(_0775_)
);

INV_X1 _1387_ (
  .A(_0769_),
  .ZN(_0771_)
);

INV_X1 _1388_ (
  .A(_0856_),
  .ZN(_0862_)
);

INV_X1 _1389_ (
  .A(_0884_),
  .ZN(_0890_)
);

INV_X1 _1390_ (
  .A(_0912_),
  .ZN(_0913_)
);

INV_X1 _1391_ (
  .A(_0950_),
  .ZN(_1204_)
);

INV_X1 _1392_ (
  .A(_0955_),
  .ZN(_0956_)
);

INV_X1 _1393_ (
  .A(_0985_),
  .ZN(_1211_)
);

INV_X1 _1394_ (
  .A(_0988_),
  .ZN(_0989_)
);

INV_X1 _1395_ (
  .A(_1026_),
  .ZN(_1028_)
);

INV_X1 _1396_ (
  .A(_1037_),
  .ZN(_1038_)
);

INV_X1 _1397_ (
  .A(_1056_),
  .ZN(_1057_)
);

INV_X1 _1398_ (
  .A(_1079_),
  .ZN(_1080_)
);

INV_X1 _1399_ (
  .A(_0689_),
  .ZN(_0699_)
);

INV_X1 _1400_ (
  .A(_0751_),
  .ZN(_0745_)
);

INV_X1 _1401_ (
  .A(_0776_),
  .ZN(_0770_)
);

INV_X1 _1402_ (
  .A(_0855_),
  .ZN(_0891_)
);

INV_X1 _1403_ (
  .A(_0883_),
  .ZN(_0924_)
);

INV_X1 _1404_ (
  .A(_0954_),
  .ZN(_0996_)
);

INV_X1 _1405_ (
  .A(_1007_),
  .ZN(_1039_)
);

INV_X1 _1406_ (
  .A(_1025_),
  .ZN(_1058_)
);

INV_X1 _1407_ (
  .A(_0702_),
  .ZN(_1141_)
);

INV_X1 _1408_ (
  .A(_0714_),
  .ZN(_0715_)
);

INV_X1 _1409_ (
  .A(_0711_),
  .ZN(_1150_)
);

INV_X1 _1410_ (
  .A(_0734_),
  .ZN(_1154_)
);

NAND2_X1 _1411_ (
  .A1(_0326_),
  .A2(_0351_),
  .ZN(_0366_)
);

INV_X1 _1412_ (
  .A(_0366_),
  .ZN(_0748_)
);

INV_X1 _1413_ (
  .A(_0723_),
  .ZN(_0774_)
);

INV_X1 _1414_ (
  .A(_0756_),
  .ZN(_0765_)
);

INV_X1 _1415_ (
  .A(_0728_),
  .ZN(_1163_)
);

INV_X1 _1416_ (
  .A(_0773_),
  .ZN(_0778_)
);

INV_X1 _1417_ (
  .A(_0789_),
  .ZN(_1171_)
);

INV_X1 _1418_ (
  .A(_0743_),
  .ZN(_0811_)
);

INV_X1 _1419_ (
  .A(_0820_),
  .ZN(_1179_)
);

INV_X1 _1420_ (
  .A(_0836_),
  .ZN(_0838_)
);

INV_X1 _1421_ (
  .A(_0809_),
  .ZN(_0837_)
);

INV_X1 _1422_ (
  .A(_0846_),
  .ZN(_0848_)
);

INV_X1 _1423_ (
  .A(_0869_),
  .ZN(_0908_)
);

INV_X1 _1424_ (
  .A(_0880_),
  .ZN(_1199_)
);

INV_X1 _1425_ (
  .A(_0946_),
  .ZN(_0947_)
);

INV_X1 _1426_ (
  .A(_0931_),
  .ZN(_0974_)
);

INV_X1 _1427_ (
  .A(_0945_),
  .ZN(_0982_)
);

INV_X1 _1428_ (
  .A(_0943_),
  .ZN(_1210_)
);

INV_X1 _1429_ (
  .A(_0991_),
  .ZN(_1216_)
);

INV_X1 _1430_ (
  .A(_0963_),
  .ZN(_1009_)
);

INV_X1 _1431_ (
  .A(_1017_),
  .ZN(_1018_)
);

INV_X1 _1432_ (
  .A(_0990_),
  .ZN(_1222_)
);

INV_X1 _1433_ (
  .A(_1046_),
  .ZN(_1047_)
);

INV_X1 _1434_ (
  .A(_1040_),
  .ZN(_1075_)
);

INV_X1 _1435_ (
  .A(_1082_),
  .ZN(_1083_)
);

INV_X1 _1436_ (
  .A(_0701_),
  .ZN(_0716_)
);

INV_X1 _1437_ (
  .A(_0762_),
  .ZN(_0766_)
);

INV_X1 _1438_ (
  .A(_0783_),
  .ZN(_0779_)
);

INV_X1 _1439_ (
  .A(_0788_),
  .ZN(_1165_)
);

INV_X1 _1440_ (
  .A(_0810_),
  .ZN(_0812_)
);

INV_X1 _1441_ (
  .A(_0761_),
  .ZN(_0813_)
);

INV_X1 _1442_ (
  .A(_0803_),
  .ZN(_0839_)
);

INV_X1 _1443_ (
  .A(_0819_),
  .ZN(_0849_)
);

INV_X1 _1444_ (
  .A(_0907_),
  .ZN(_0909_)
);

INV_X1 _1445_ (
  .A(_0914_),
  .ZN(_0948_)
);

INV_X1 _1446_ (
  .A(_0917_),
  .ZN(_1205_)
);

INV_X1 _1447_ (
  .A(_0935_),
  .ZN(_0973_)
);

INV_X1 _1448_ (
  .A(_0972_),
  .ZN(_0975_)
);

INV_X1 _1449_ (
  .A(_0939_),
  .ZN(_0976_)
);

INV_X1 _1450_ (
  .A(_0980_),
  .ZN(_0983_)
);

INV_X1 _1451_ (
  .A(_0967_),
  .ZN(_1006_)
);

INV_X1 _1452_ (
  .A(_0971_),
  .ZN(_1010_)
);

INV_X1 _1453_ (
  .A(_0902_),
  .ZN(_0942_)
);

INV_X1 _1454_ (
  .A(_1016_),
  .ZN(_1048_)
);

INV_X1 _1455_ (
  .A(_1045_),
  .ZN(_1084_)
);

INV_X1 _1456_ (
  .A(_1153_),
  .ZN(_0732_)
);

INV_X1 _1457_ (
  .A(_1170_),
  .ZN(_0790_)
);

INV_X1 _1458_ (
  .A(_1178_),
  .ZN(_0818_)
);

INV_X1 _1459_ (
  .A(_1187_),
  .ZN(_0844_)
);

INV_X1 _1460_ (
  .A(_1194_),
  .ZN(_0876_)
);

INV_X1 _1461_ (
  .A(_1219_),
  .ZN(_1015_)
);

INV_X1 _1462_ (
  .A(_1228_),
  .ZN(_1044_)
);

INV_X1 _1463_ (
  .A(_1140_),
  .ZN(_0700_)
);

INV_X1 _1464_ (
  .A(_1164_),
  .ZN(_0784_)
);

INV_X1 _1465_ (
  .A(_0941_),
  .ZN(_0937_)
);

INV_X1 _1466_ (
  .A(_1173_),
  .ZN(_0791_)
);

BUF_X1 _1467_ (
  .A(ena),
  .Z(_0367_)
);

BUF_X1 _1468_ (
  .A(_0367_),
  .Z(_0368_)
);

NAND3_X1 _1469_ (
  .A1(din[0]),
  .A2(_0329_),
  .A3(_0368_),
  .ZN(_0369_)
);

INV_X1 _1470_ (
  .A(\ext_mult_res[0] ),
  .ZN(_0370_)
);

BUF_X1 _1471_ (
  .A(_0367_),
  .Z(_0371_)
);

BUF_X1 _1472_ (
  .A(_0371_),
  .Z(_0372_)
);

OAI21_X1 _1473_ (
  .A(_0369_),
  .B1(_0370_),
  .B2(_0372_),
  .ZN(_0000_)
);

BUF_X1 _1474_ (
  .A(_0367_),
  .Z(_0373_)
);

MUX2_X1 _1475_ (
  .A(\ext_mult_res[1] ),
  .B(_1133_),
  .S(_0373_),
  .Z(_0001_)
);

BUF_X4 _1476_ (
  .A(_0371_),
  .Z(_0374_)
);

NAND2_X1 _1477_ (
  .A1(_0374_),
  .A2(_1135_),
  .ZN(_0375_)
);

INV_X1 _1478_ (
  .A(\ext_mult_res[2] ),
  .ZN(_0376_)
);

OAI21_X1 _1479_ (
  .A(_0375_),
  .B1(_0376_),
  .B2(_0372_),
  .ZN(_0002_)
);

NAND2_X1 _1480_ (
  .A1(_0374_),
  .A2(_1137_),
  .ZN(_0377_)
);

INV_X1 _1481_ (
  .A(\ext_mult_res[3] ),
  .ZN(_0378_)
);

OAI21_X1 _1482_ (
  .A(_0377_),
  .B1(_0378_),
  .B2(_0372_),
  .ZN(_0003_)
);

NAND2_X1 _1483_ (
  .A1(_0374_),
  .A2(_1145_),
  .ZN(_0379_)
);

INV_X1 _1484_ (
  .A(\ext_mult_res[4] ),
  .ZN(_0380_)
);

OAI21_X1 _1485_ (
  .A(_0379_),
  .B1(_0380_),
  .B2(_0372_),
  .ZN(_0004_)
);

MUX2_X1 _1486_ (
  .A(\ext_mult_res[5] ),
  .B(_1149_),
  .S(_0373_),
  .Z(_0005_)
);

NAND2_X1 _1487_ (
  .A1(_0372_),
  .A2(_1160_),
  .ZN(_0381_)
);

INV_X1 _1488_ (
  .A(\ext_mult_res[6] ),
  .ZN(_0382_)
);

OAI21_X1 _1489_ (
  .A(_0381_),
  .B1(_0382_),
  .B2(_0372_),
  .ZN(_0006_)
);

NAND2_X1 _1490_ (
  .A1(_0374_),
  .A2(_1234_),
  .ZN(_0383_)
);

INV_X1 _1491_ (
  .A(\ext_mult_res[7] ),
  .ZN(_0384_)
);

OAI21_X1 _1492_ (
  .A(_0383_),
  .B1(_0384_),
  .B2(_0372_),
  .ZN(_0007_)
);

INV_X1 _1493_ (
  .A(_0367_),
  .ZN(_0385_)
);

NAND2_X1 _1494_ (
  .A1(_0385_),
  .A2(\ext_mult_res[8] ),
  .ZN(_0386_)
);

BUF_X1 _1495_ (
  .A(_0385_),
  .Z(_0387_)
);

OAI21_X1 _1496_ (
  .A(_0386_),
  .B1(_0794_),
  .B2(_0387_),
  .ZN(_0008_)
);

INV_X1 _1497_ (
  .A(_0793_),
  .ZN(_0388_)
);

NAND2_X1 _1498_ (
  .A1(_0388_),
  .A2(_1185_),
  .ZN(_0389_)
);

INV_X1 _1499_ (
  .A(_1185_),
  .ZN(_0390_)
);

NAND2_X1 _1500_ (
  .A1(_0390_),
  .A2(_0793_),
  .ZN(_0391_)
);

NAND3_X1 _1501_ (
  .A1(_0389_),
  .A2(_0391_),
  .A3(_0374_),
  .ZN(_0392_)
);

INV_X1 _1502_ (
  .A(\ext_mult_res[9] ),
  .ZN(_0393_)
);

OAI21_X1 _1503_ (
  .A(_0392_),
  .B1(_0393_),
  .B2(_0372_),
  .ZN(_0009_)
);

NOR2_X1 _1504_ (
  .A1(\ext_mult_res[10] ),
  .A2(_0373_),
  .ZN(_0394_)
);

INV_X1 _1505_ (
  .A(_1184_),
  .ZN(_0395_)
);

INV_X1 _1506_ (
  .A(_1174_),
  .ZN(_0396_)
);

OAI21_X1 _1507_ (
  .A(_0395_),
  .B1(_0390_),
  .B2(_0396_),
  .ZN(_0397_)
);

INV_X1 _1508_ (
  .A(_0397_),
  .ZN(_0398_)
);

NAND2_X1 _1509_ (
  .A1(_1185_),
  .A2(_1175_),
  .ZN(_0399_)
);

OAI21_X1 _1510_ (
  .A(_0398_),
  .B1(_0792_),
  .B2(_0399_),
  .ZN(_0400_)
);

BUF_X1 _1511_ (
  .A(_1191_),
  .Z(_0401_)
);

XNOR2_X1 _1512_ (
  .A(_0400_),
  .B(_0401_),
  .ZN(_0402_)
);

BUF_X1 _1513_ (
  .A(_0371_),
  .Z(_0403_)
);

AOI21_X1 _1514_ (
  .A(_0394_),
  .B1(_0402_),
  .B2(_0403_),
  .ZN(_0010_)
);

NOR2_X1 _1515_ (
  .A1(\ext_mult_res[11] ),
  .A2(_0373_),
  .ZN(_0404_)
);

INV_X1 _1516_ (
  .A(_1190_),
  .ZN(_0405_)
);

INV_X1 _1517_ (
  .A(_0401_),
  .ZN(_0406_)
);

OAI21_X1 _1518_ (
  .A(_0405_),
  .B1(_0406_),
  .B2(_0395_),
  .ZN(_0407_)
);

NAND2_X1 _1519_ (
  .A1(_1185_),
  .A2(_0401_),
  .ZN(_0408_)
);

INV_X1 _1520_ (
  .A(_0408_),
  .ZN(_0409_)
);

AOI21_X1 _1521_ (
  .A(_0407_),
  .B1(_0409_),
  .B2(_0388_),
  .ZN(_0410_)
);

INV_X1 _1522_ (
  .A(_1198_),
  .ZN(_0411_)
);

XNOR2_X1 _1523_ (
  .A(_0410_),
  .B(_0411_),
  .ZN(_0412_)
);

AOI21_X1 _1524_ (
  .A(_0404_),
  .B1(_0412_),
  .B2(_0403_),
  .ZN(_0011_)
);

NOR2_X1 _1525_ (
  .A1(\ext_mult_res[12] ),
  .A2(_0373_),
  .ZN(_0413_)
);

INV_X1 _1526_ (
  .A(_1197_),
  .ZN(_0414_)
);

OAI21_X1 _1527_ (
  .A(_0414_),
  .B1(_0411_),
  .B2(_0405_),
  .ZN(_0415_)
);

INV_X1 _1528_ (
  .A(_0415_),
  .ZN(_0416_)
);

NAND2_X1 _1529_ (
  .A1(_0401_),
  .A2(_1198_),
  .ZN(_0417_)
);

OAI21_X1 _1530_ (
  .A(_0416_),
  .B1(_0398_),
  .B2(_0417_),
  .ZN(_0418_)
);

NOR2_X1 _1531_ (
  .A1(_0399_),
  .A2(_0417_),
  .ZN(_0419_)
);

AOI21_X1 _1532_ (
  .A(_0418_),
  .B1(_0419_),
  .B2(_1177_),
  .ZN(_0420_)
);

INV_X1 _1533_ (
  .A(_1203_),
  .ZN(_0421_)
);

XNOR2_X1 _1534_ (
  .A(_0420_),
  .B(_0421_),
  .ZN(_0422_)
);

AOI21_X1 _1535_ (
  .A(_0413_),
  .B1(_0422_),
  .B2(_0403_),
  .ZN(_0012_)
);

NOR2_X1 _1536_ (
  .A1(\ext_mult_res[13] ),
  .A2(_0373_),
  .ZN(_0423_)
);

INV_X1 _1537_ (
  .A(_1202_),
  .ZN(_0424_)
);

OAI21_X1 _1538_ (
  .A(_0424_),
  .B1(_0421_),
  .B2(_0414_),
  .ZN(_0425_)
);

INV_X1 _1539_ (
  .A(_0425_),
  .ZN(_0426_)
);

INV_X1 _1540_ (
  .A(_0407_),
  .ZN(_0427_)
);

NAND2_X1 _1541_ (
  .A1(_1198_),
  .A2(_1203_),
  .ZN(_0428_)
);

OAI21_X1 _1542_ (
  .A(_0426_),
  .B1(_0427_),
  .B2(_0428_),
  .ZN(_0429_)
);

NOR2_X1 _1543_ (
  .A1(_0408_),
  .A2(_0428_),
  .ZN(_0430_)
);

AOI21_X1 _1544_ (
  .A(_0429_),
  .B1(_0430_),
  .B2(_0388_),
  .ZN(_0431_)
);

INV_X1 _1545_ (
  .A(_1209_),
  .ZN(_0432_)
);

XNOR2_X1 _1546_ (
  .A(_0431_),
  .B(_0432_),
  .ZN(_0433_)
);

AOI21_X1 _1547_ (
  .A(_0423_),
  .B1(_0433_),
  .B2(_0403_),
  .ZN(_0013_)
);

NOR2_X1 _1548_ (
  .A1(\ext_mult_res[14] ),
  .A2(_0373_),
  .ZN(_0434_)
);

INV_X1 _1549_ (
  .A(_1208_),
  .ZN(_0435_)
);

OAI21_X1 _1550_ (
  .A(_0435_),
  .B1(_0432_),
  .B2(_0424_),
  .ZN(_0436_)
);

INV_X1 _1551_ (
  .A(_0436_),
  .ZN(_0437_)
);

NAND2_X1 _1552_ (
  .A1(_1203_),
  .A2(_1209_),
  .ZN(_0438_)
);

OAI21_X1 _1553_ (
  .A(_0437_),
  .B1(_0416_),
  .B2(_0438_),
  .ZN(_0439_)
);

NOR2_X1 _1554_ (
  .A1(_0417_),
  .A2(_0438_),
  .ZN(_0440_)
);

AOI21_X1 _1555_ (
  .A(_0439_),
  .B1(_0440_),
  .B2(_0400_),
  .ZN(_0441_)
);

INV_X1 _1556_ (
  .A(_1215_),
  .ZN(_0442_)
);

XNOR2_X1 _1557_ (
  .A(_0441_),
  .B(_0442_),
  .ZN(_0443_)
);

AOI21_X1 _1558_ (
  .A(_0434_),
  .B1(_0443_),
  .B2(_0403_),
  .ZN(_0014_)
);

NAND2_X1 _1559_ (
  .A1(_1209_),
  .A2(_1215_),
  .ZN(_0444_)
);

NOR3_X1 _1560_ (
  .A1(_0410_),
  .A2(_0428_),
  .A3(_0444_),
  .ZN(_0445_)
);

INV_X1 _1561_ (
  .A(_1214_),
  .ZN(_0446_)
);

OAI21_X1 _1562_ (
  .A(_0446_),
  .B1(_0442_),
  .B2(_0435_),
  .ZN(_0447_)
);

INV_X1 _1563_ (
  .A(_0447_),
  .ZN(_0448_)
);

OAI21_X1 _1564_ (
  .A(_0448_),
  .B1(_0426_),
  .B2(_0444_),
  .ZN(_0449_)
);

OR2_X1 _1565_ (
  .A1(_0445_),
  .A2(_0449_),
  .ZN(_0450_)
);

BUF_X1 _1566_ (
  .A(_1221_),
  .Z(_0451_)
);

OR2_X1 _1567_ (
  .A1(_0450_),
  .A2(_0451_),
  .ZN(_0452_)
);

NAND2_X1 _1568_ (
  .A1(_0450_),
  .A2(_0451_),
  .ZN(_0453_)
);

NAND3_X1 _1569_ (
  .A1(_0452_),
  .A2(_0374_),
  .A3(_0453_),
  .ZN(_0454_)
);

INV_X1 _1570_ (
  .A(\ext_mult_res[15] ),
  .ZN(_0455_)
);

OAI21_X1 _1571_ (
  .A(_0454_),
  .B1(_0455_),
  .B2(_0372_),
  .ZN(_0015_)
);

NOR2_X1 _1572_ (
  .A1(\ext_mult_res[16] ),
  .A2(_0373_),
  .ZN(_0456_)
);

INV_X1 _1573_ (
  .A(_1220_),
  .ZN(_0457_)
);

INV_X1 _1574_ (
  .A(_0451_),
  .ZN(_0458_)
);

OAI21_X1 _1575_ (
  .A(_0457_),
  .B1(_0458_),
  .B2(_0446_),
  .ZN(_0459_)
);

INV_X1 _1576_ (
  .A(_0459_),
  .ZN(_0460_)
);

NAND2_X1 _1577_ (
  .A1(_1215_),
  .A2(_0451_),
  .ZN(_0461_)
);

OAI21_X1 _1578_ (
  .A(_0460_),
  .B1(_0437_),
  .B2(_0461_),
  .ZN(_0462_)
);

NOR2_X1 _1579_ (
  .A1(_0438_),
  .A2(_0461_),
  .ZN(_0463_)
);

AOI21_X1 _1580_ (
  .A(_0462_),
  .B1(_0463_),
  .B2(_0418_),
  .ZN(_0464_)
);

NAND3_X1 _1581_ (
  .A1(_0419_),
  .A2(_0463_),
  .A3(_1177_),
  .ZN(_0465_)
);

NAND2_X1 _1582_ (
  .A1(_0464_),
  .A2(_0465_),
  .ZN(_0466_)
);

BUF_X1 _1583_ (
  .A(_1230_),
  .Z(_0467_)
);

XNOR2_X1 _1584_ (
  .A(_0466_),
  .B(_0467_),
  .ZN(_0468_)
);

AOI21_X1 _1585_ (
  .A(_0456_),
  .B1(_0468_),
  .B2(_0403_),
  .ZN(_0016_)
);

NOR2_X1 _1586_ (
  .A1(\ext_mult_res[17] ),
  .A2(_0373_),
  .ZN(_0469_)
);

INV_X1 _1587_ (
  .A(_1229_),
  .ZN(_0470_)
);

INV_X1 _1588_ (
  .A(_0467_),
  .ZN(_0471_)
);

NAND2_X1 _1589_ (
  .A1(_0451_),
  .A2(_0467_),
  .ZN(_0472_)
);

OAI221_X1 _1590_ (
  .A(_0470_),
  .B1(_0457_),
  .B2(_0471_),
  .C1(_0448_),
  .C2(_0472_),
  .ZN(_0473_)
);

INV_X1 _1591_ (
  .A(_0473_),
  .ZN(_0474_)
);

NOR2_X1 _1592_ (
  .A1(_0444_),
  .A2(_0472_),
  .ZN(_0475_)
);

NAND2_X1 _1593_ (
  .A1(_0429_),
  .A2(_0475_),
  .ZN(_0476_)
);

NAND3_X1 _1594_ (
  .A1(_0430_),
  .A2(_0475_),
  .A3(_0388_),
  .ZN(_0477_)
);

NAND3_X1 _1595_ (
  .A1(_0474_),
  .A2(_0476_),
  .A3(_0477_),
  .ZN(_0478_)
);

BUF_X1 _1596_ (
  .A(_1233_),
  .Z(_0479_)
);

XNOR2_X1 _1597_ (
  .A(_0478_),
  .B(_0479_),
  .ZN(_0480_)
);

AOI21_X1 _1598_ (
  .A(_0469_),
  .B1(_0480_),
  .B2(_0403_),
  .ZN(_0017_)
);

INV_X1 _1599_ (
  .A(_1061_),
  .ZN(_0481_)
);

INV_X1 _1600_ (
  .A(_1070_),
  .ZN(_0482_)
);

NAND2_X1 _1601_ (
  .A1(_0481_),
  .A2(_0482_),
  .ZN(_0483_)
);

NAND2_X1 _1602_ (
  .A1(_1061_),
  .A2(_1070_),
  .ZN(_0484_)
);

NAND2_X1 _1603_ (
  .A1(_0483_),
  .A2(_0484_),
  .ZN(_0485_)
);

INV_X1 _1604_ (
  .A(_0485_),
  .ZN(_0486_)
);

INV_X1 _1605_ (
  .A(_1081_),
  .ZN(_0487_)
);

NAND2_X1 _1606_ (
  .A1(_0487_),
  .A2(_1055_),
  .ZN(_0488_)
);

INV_X1 _1607_ (
  .A(_1055_),
  .ZN(_0489_)
);

NAND2_X1 _1608_ (
  .A1(_0489_),
  .A2(_1081_),
  .ZN(_0490_)
);

NAND2_X1 _1609_ (
  .A1(_0488_),
  .A2(_0490_),
  .ZN(_0491_)
);

NAND2_X1 _1610_ (
  .A1(_0486_),
  .A2(_0491_),
  .ZN(_0492_)
);

XNOR2_X1 _1611_ (
  .A(_1081_),
  .B(_1055_),
  .ZN(_0493_)
);

NAND2_X1 _1612_ (
  .A1(_0493_),
  .A2(_0485_),
  .ZN(_0494_)
);

NAND2_X1 _1613_ (
  .A1(_0492_),
  .A2(_0494_),
  .ZN(_0495_)
);

INV_X1 _1614_ (
  .A(_1224_),
  .ZN(_0496_)
);

NAND2_X1 _1615_ (
  .A1(_0496_),
  .A2(_1027_),
  .ZN(_0497_)
);

NAND2_X1 _1616_ (
  .A1(_1224_),
  .A2(_0987_),
  .ZN(_0498_)
);

NAND2_X1 _1617_ (
  .A1(_0497_),
  .A2(_0498_),
  .ZN(_0499_)
);

NAND2_X1 _1618_ (
  .A1(_0499_),
  .A2(_1023_),
  .ZN(_0500_)
);

NAND3_X1 _1619_ (
  .A1(_0497_),
  .A2(_1052_),
  .A3(_0498_),
  .ZN(_0501_)
);

NAND2_X2 _1620_ (
  .A1(_0500_),
  .A2(_0501_),
  .ZN(_0502_)
);

XNOR2_X1 _1621_ (
  .A(_0495_),
  .B(_0502_),
  .ZN(_0503_)
);

INV_X1 _1622_ (
  .A(_1005_),
  .ZN(_0504_)
);

XNOR2_X1 _1623_ (
  .A(_0504_),
  .B(_1059_),
  .ZN(_0505_)
);

XNOR2_X1 _1624_ (
  .A(_1063_),
  .B(_1065_),
  .ZN(_0506_)
);

NAND2_X1 _1625_ (
  .A1(_0505_),
  .A2(_0506_),
  .ZN(_0507_)
);

NAND2_X1 _1626_ (
  .A1(_1063_),
  .A2(_1065_),
  .ZN(_0508_)
);

INV_X1 _1627_ (
  .A(_0508_),
  .ZN(_0509_)
);

NOR2_X1 _1628_ (
  .A1(_1063_),
  .A2(_1065_),
  .ZN(_0510_)
);

NOR2_X1 _1629_ (
  .A1(_0509_),
  .A2(_0510_),
  .ZN(_0511_)
);

XNOR2_X1 _1630_ (
  .A(_1005_),
  .B(_1059_),
  .ZN(_0512_)
);

NAND2_X1 _1631_ (
  .A1(_0511_),
  .A2(_0512_),
  .ZN(_0513_)
);

NAND2_X1 _1632_ (
  .A1(_0507_),
  .A2(_0513_),
  .ZN(_0514_)
);

INV_X1 _1633_ (
  .A(_0514_),
  .ZN(_0515_)
);

NAND2_X4 _1634_ (
  .A1(_0960_),
  .A2(_0993_),
  .ZN(_0516_)
);

NAND3_X4 _1635_ (
  .A1(_0350_),
  .A2(_0351_),
  .A3(_0356_),
  .ZN(_0517_)
);

NAND2_X4 _1636_ (
  .A1(_0516_),
  .A2(_0517_),
  .ZN(_0518_)
);

NAND2_X2 _1637_ (
  .A1(_0518_),
  .A2(_1053_),
  .ZN(_0519_)
);

NAND3_X1 _1638_ (
  .A1(_0516_),
  .A2(_0517_),
  .A3(_0358_),
  .ZN(_0520_)
);

NAND2_X2 _1639_ (
  .A1(_0519_),
  .A2(_0520_),
  .ZN(_0521_)
);

NAND2_X1 _1640_ (
  .A1(_0515_),
  .A2(_0521_),
  .ZN(_0522_)
);

NAND2_X2 _1641_ (
  .A1(_0518_),
  .A2(_1024_),
  .ZN(_0523_)
);

INV_X1 _1642_ (
  .A(_0358_),
  .ZN(_0524_)
);

NAND3_X1 _1643_ (
  .A1(_0516_),
  .A2(_0517_),
  .A3(_0524_),
  .ZN(_0525_)
);

NAND2_X2 _1644_ (
  .A1(_0523_),
  .A2(_0525_),
  .ZN(_0526_)
);

NAND2_X1 _1645_ (
  .A1(_0526_),
  .A2(_0514_),
  .ZN(_0527_)
);

NAND2_X2 _1646_ (
  .A1(_0522_),
  .A2(_0527_),
  .ZN(_0528_)
);

NAND2_X1 _1647_ (
  .A1(_0503_),
  .A2(_0528_),
  .ZN(_0529_)
);

NAND2_X1 _1648_ (
  .A1(_0515_),
  .A2(_0526_),
  .ZN(_0530_)
);

NAND2_X1 _1649_ (
  .A1(_0521_),
  .A2(_0514_),
  .ZN(_0531_)
);

NAND2_X2 _1650_ (
  .A1(_0530_),
  .A2(_0531_),
  .ZN(_0532_)
);

XNOR2_X1 _1651_ (
  .A(_0491_),
  .B(_0485_),
  .ZN(_0533_)
);

NAND2_X1 _1652_ (
  .A1(_0533_),
  .A2(_0502_),
  .ZN(_0534_)
);

INV_X1 _1653_ (
  .A(_0502_),
  .ZN(_0535_)
);

NAND2_X1 _1654_ (
  .A1(_0495_),
  .A2(_0535_),
  .ZN(_0536_)
);

NAND2_X1 _1655_ (
  .A1(_0534_),
  .A2(_0536_),
  .ZN(_0537_)
);

NAND2_X1 _1656_ (
  .A1(_0532_),
  .A2(_0537_),
  .ZN(_0538_)
);

NAND2_X1 _1657_ (
  .A1(_0529_),
  .A2(_0538_),
  .ZN(_0539_)
);

OR2_X1 _1658_ (
  .A1(_1086_),
  .A2(_1078_),
  .ZN(_0540_)
);

NAND2_X1 _1659_ (
  .A1(_1078_),
  .A2(_1086_),
  .ZN(_0541_)
);

NAND2_X1 _1660_ (
  .A1(_0540_),
  .A2(_0541_),
  .ZN(_0542_)
);

NAND2_X4 _1661_ (
  .A1(_0542_),
  .A2(_0764_),
  .ZN(_0543_)
);

NAND3_X2 _1662_ (
  .A1(_0540_),
  .A2(_0760_),
  .A3(_0541_),
  .ZN(_0544_)
);

NAND2_X2 _1663_ (
  .A1(_0543_),
  .A2(_0544_),
  .ZN(_0545_)
);

XOR2_X1 _1664_ (
  .A(_1068_),
  .B(_1231_),
  .Z(_0546_)
);

INV_X1 _1665_ (
  .A(_0546_),
  .ZN(_0547_)
);

NAND2_X2 _1666_ (
  .A1(_0545_),
  .A2(_0547_),
  .ZN(_0548_)
);

NAND3_X2 _1667_ (
  .A1(_0543_),
  .A2(_0544_),
  .A3(_0546_),
  .ZN(_0549_)
);

NAND2_X2 _1668_ (
  .A1(_0548_),
  .A2(_0549_),
  .ZN(_0550_)
);

XNOR2_X1 _1669_ (
  .A(_0967_),
  .B(_0903_),
  .ZN(_0551_)
);

XNOR2_X1 _1670_ (
  .A(_0874_),
  .B(_1073_),
  .ZN(_0552_)
);

XNOR2_X1 _1671_ (
  .A(_0551_),
  .B(_0552_),
  .ZN(_0553_)
);

INV_X1 _1672_ (
  .A(_0553_),
  .ZN(_0554_)
);

NAND2_X2 _1673_ (
  .A1(_0550_),
  .A2(_0554_),
  .ZN(_0555_)
);

NAND3_X1 _1674_ (
  .A1(_0548_),
  .A2(_0549_),
  .A3(_0553_),
  .ZN(_0556_)
);

NAND2_X2 _1675_ (
  .A1(_0555_),
  .A2(_0556_),
  .ZN(_0557_)
);

INV_X1 _1676_ (
  .A(_0557_),
  .ZN(_0558_)
);

NAND2_X2 _1677_ (
  .A1(_0539_),
  .A2(_0558_),
  .ZN(_0559_)
);

NAND2_X1 _1678_ (
  .A1(_0503_),
  .A2(_0532_),
  .ZN(_0560_)
);

NAND2_X1 _1679_ (
  .A1(_0528_),
  .A2(_0537_),
  .ZN(_0561_)
);

NAND2_X2 _1680_ (
  .A1(_0560_),
  .A2(_0561_),
  .ZN(_0562_)
);

NAND2_X2 _1681_ (
  .A1(_0562_),
  .A2(_0557_),
  .ZN(_0563_)
);

NAND2_X2 _1682_ (
  .A1(_0559_),
  .A2(_0563_),
  .ZN(_0564_)
);

INV_X1 _1683_ (
  .A(_0479_),
  .ZN(_0565_)
);

NOR3_X1 _1684_ (
  .A1(_0461_),
  .A2(_0471_),
  .A3(_0565_),
  .ZN(_0566_)
);

NAND3_X1 _1685_ (
  .A1(_0400_),
  .A2(_0440_),
  .A3(_0566_),
  .ZN(_0567_)
);

NAND3_X1 _1686_ (
  .A1(_0459_),
  .A2(_0467_),
  .A3(_0479_),
  .ZN(_0568_)
);

INV_X1 _1687_ (
  .A(_1232_),
  .ZN(_0569_)
);

NAND2_X1 _1688_ (
  .A1(_0479_),
  .A2(_1229_),
  .ZN(_0570_)
);

NAND3_X1 _1689_ (
  .A1(_0568_),
  .A2(_0569_),
  .A3(_0570_),
  .ZN(_0571_)
);

INV_X1 _1690_ (
  .A(_0571_),
  .ZN(_0572_)
);

NAND2_X1 _1691_ (
  .A1(_0439_),
  .A2(_0566_),
  .ZN(_0573_)
);

AND3_X1 _1692_ (
  .A1(_0567_),
  .A2(_0572_),
  .A3(_0573_),
  .ZN(_0574_)
);

INV_X1 _1693_ (
  .A(_0574_),
  .ZN(_0575_)
);

NAND2_X2 _1694_ (
  .A1(_0564_),
  .A2(_0575_),
  .ZN(_0576_)
);

NAND3_X1 _1695_ (
  .A1(_0559_),
  .A2(_0563_),
  .A3(_0574_),
  .ZN(_0577_)
);

NAND3_X1 _1696_ (
  .A1(_0576_),
  .A2(_0577_),
  .A3(_0374_),
  .ZN(_0578_)
);

NAND2_X1 _1697_ (
  .A1(_0387_),
  .A2(\ext_mult_res[18] ),
  .ZN(_0579_)
);

NAND2_X1 _1698_ (
  .A1(_0578_),
  .A2(_0579_),
  .ZN(_0018_)
);

NAND2_X1 _1699_ (
  .A1(_0385_),
  .A2(result[0]),
  .ZN(_0580_)
);

BUF_X1 _1700_ (
  .A(dclr),
  .Z(_0581_)
);

OAI21_X1 _1701_ (
  .A(_0368_),
  .B1(_1089_),
  .B2(_0581_),
  .ZN(_0582_)
);

INV_X1 _1702_ (
  .A(_0581_),
  .ZN(_0583_)
);

BUF_X1 _1703_ (
  .A(_0583_),
  .Z(_0584_)
);

NOR2_X1 _1704_ (
  .A1(_0584_),
  .A2(\ext_mult_res[0] ),
  .ZN(_0585_)
);

OAI21_X1 _1705_ (
  .A(_0580_),
  .B1(_0582_),
  .B2(_0585_),
  .ZN(_0019_)
);

NAND2_X1 _1706_ (
  .A1(_0385_),
  .A2(result[1]),
  .ZN(_0586_)
);

OAI21_X1 _1707_ (
  .A(_0368_),
  .B1(_0581_),
  .B2(_0680_),
  .ZN(_0587_)
);

NOR2_X1 _1708_ (
  .A1(_0584_),
  .A2(\ext_mult_res[1] ),
  .ZN(_0588_)
);

OAI21_X1 _1709_ (
  .A(_0586_),
  .B1(_0587_),
  .B2(_0588_),
  .ZN(_0020_)
);

INV_X1 _1710_ (
  .A(_1093_),
  .ZN(_0589_)
);

NOR2_X1 _1711_ (
  .A1(_0589_),
  .A2(_0679_),
  .ZN(_0590_)
);

INV_X1 _1712_ (
  .A(_0590_),
  .ZN(_0591_)
);

NAND2_X1 _1713_ (
  .A1(_0589_),
  .A2(_0679_),
  .ZN(_0592_)
);

NAND3_X1 _1714_ (
  .A1(_0591_),
  .A2(_0583_),
  .A3(_0592_),
  .ZN(_0593_)
);

BUF_X2 _1715_ (
  .A(_0583_),
  .Z(_0594_)
);

OAI21_X1 _1716_ (
  .A(_0593_),
  .B1(_0594_),
  .B2(_0376_),
  .ZN(_0595_)
);

MUX2_X1 _1717_ (
  .A(result[2]),
  .B(_0595_),
  .S(_0373_),
  .Z(_0021_)
);

OAI21_X1 _1718_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(_0378_),
  .ZN(_0596_)
);

NAND2_X1 _1719_ (
  .A1(_1088_),
  .A2(_1091_),
  .ZN(_0597_)
);

INV_X1 _1720_ (
  .A(_1090_),
  .ZN(_0598_)
);

INV_X1 _1721_ (
  .A(_1092_),
  .ZN(_0599_)
);

NAND3_X1 _1722_ (
  .A1(_0597_),
  .A2(_0598_),
  .A3(_0599_),
  .ZN(_0600_)
);

NAND2_X1 _1723_ (
  .A1(_0589_),
  .A2(_0599_),
  .ZN(_0601_)
);

NAND2_X1 _1724_ (
  .A1(_0600_),
  .A2(_0601_),
  .ZN(_0602_)
);

XNOR2_X1 _1725_ (
  .A(_0602_),
  .B(_1095_),
  .ZN(_0603_)
);

BUF_X1 _1726_ (
  .A(_0583_),
  .Z(_0604_)
);

AOI21_X1 _1727_ (
  .A(_0596_),
  .B1(_0603_),
  .B2(_0604_),
  .ZN(_0605_)
);

INV_X1 _1728_ (
  .A(result[3]),
  .ZN(_0606_)
);

AOI21_X1 _1729_ (
  .A(_0605_),
  .B1(_0606_),
  .B2(_0387_),
  .ZN(_0022_)
);

OAI21_X1 _1730_ (
  .A(_0367_),
  .B1(_0583_),
  .B2(_0380_),
  .ZN(_0607_)
);

INV_X1 _1731_ (
  .A(_1094_),
  .ZN(_0608_)
);

INV_X1 _1732_ (
  .A(_1095_),
  .ZN(_0609_)
);

OAI21_X1 _1733_ (
  .A(_0608_),
  .B1(_0609_),
  .B2(_0599_),
  .ZN(_0610_)
);

INV_X1 _1734_ (
  .A(_0610_),
  .ZN(_0611_)
);

OAI21_X4 _1735_ (
  .A(_0611_),
  .B1(_0609_),
  .B2(_0591_),
  .ZN(_0612_)
);

INV_X1 _1736_ (
  .A(_1097_),
  .ZN(_0613_)
);

XNOR2_X1 _1737_ (
  .A(_0612_),
  .B(_0613_),
  .ZN(_0614_)
);

AOI21_X1 _1738_ (
  .A(_0607_),
  .B1(_0614_),
  .B2(_0604_),
  .ZN(_0615_)
);

INV_X1 _1739_ (
  .A(result[4]),
  .ZN(_0616_)
);

AOI21_X1 _1740_ (
  .A(_0615_),
  .B1(_0616_),
  .B2(_0387_),
  .ZN(_0023_)
);

NAND2_X1 _1741_ (
  .A1(_1095_),
  .A2(_1097_),
  .ZN(_0617_)
);

INV_X1 _1742_ (
  .A(_0617_),
  .ZN(_0618_)
);

NAND3_X1 _1743_ (
  .A1(_0600_),
  .A2(_0601_),
  .A3(_0618_),
  .ZN(_0619_)
);

INV_X1 _1744_ (
  .A(_1096_),
  .ZN(_0620_)
);

OAI21_X1 _1745_ (
  .A(_0620_),
  .B1(_0613_),
  .B2(_0608_),
  .ZN(_0621_)
);

INV_X1 _1746_ (
  .A(_0621_),
  .ZN(_0622_)
);

NAND2_X1 _1747_ (
  .A1(_0619_),
  .A2(_0622_),
  .ZN(_0623_)
);

BUF_X2 _1748_ (
  .A(_1099_),
  .Z(_0624_)
);

XNOR2_X1 _1749_ (
  .A(_0623_),
  .B(_0624_),
  .ZN(_0625_)
);

AOI21_X1 _1750_ (
  .A(_0385_),
  .B1(_0625_),
  .B2(_0594_),
  .ZN(_0626_)
);

OAI21_X1 _1751_ (
  .A(_0626_),
  .B1(_0584_),
  .B2(\ext_mult_res[5] ),
  .ZN(_0627_)
);

INV_X1 _1752_ (
  .A(result[5]),
  .ZN(_0628_)
);

OAI21_X1 _1753_ (
  .A(_0627_),
  .B1(_0403_),
  .B2(_0628_),
  .ZN(_0024_)
);

INV_X1 _1754_ (
  .A(_1098_),
  .ZN(_0629_)
);

INV_X1 _1755_ (
  .A(_0624_),
  .ZN(_0630_)
);

OAI21_X1 _1756_ (
  .A(_0629_),
  .B1(_0630_),
  .B2(_0620_),
  .ZN(_0631_)
);

INV_X1 _1757_ (
  .A(_0631_),
  .ZN(_0632_)
);

INV_X1 _1758_ (
  .A(_0612_),
  .ZN(_0633_)
);

NAND2_X1 _1759_ (
  .A1(_1097_),
  .A2(_0624_),
  .ZN(_0634_)
);

OAI21_X1 _1760_ (
  .A(_0632_),
  .B1(_0633_),
  .B2(_0634_),
  .ZN(_0635_)
);

CLKBUF_X2 _1761_ (
  .A(_1101_),
  .Z(_0636_)
);

XNOR2_X1 _1762_ (
  .A(_0635_),
  .B(_0636_),
  .ZN(_0041_)
);

NAND2_X1 _1763_ (
  .A1(_0041_),
  .A2(_0604_),
  .ZN(_0042_)
);

NAND2_X1 _1764_ (
  .A1(_0382_),
  .A2(_0581_),
  .ZN(_0043_)
);

NAND3_X1 _1765_ (
  .A1(_0042_),
  .A2(_0374_),
  .A3(_0043_),
  .ZN(_0044_)
);

INV_X1 _1766_ (
  .A(result[6]),
  .ZN(_0045_)
);

OAI21_X1 _1767_ (
  .A(_0044_),
  .B1(_0403_),
  .B2(_0045_),
  .ZN(_0025_)
);

NAND2_X1 _1768_ (
  .A1(_0636_),
  .A2(_1098_),
  .ZN(_0046_)
);

INV_X1 _1769_ (
  .A(_1100_),
  .ZN(_0047_)
);

NAND2_X1 _1770_ (
  .A1(_0046_),
  .A2(_0047_),
  .ZN(_0048_)
);

INV_X1 _1771_ (
  .A(_0048_),
  .ZN(_0049_)
);

NAND2_X1 _1772_ (
  .A1(_0624_),
  .A2(_0636_),
  .ZN(_0050_)
);

OAI21_X1 _1773_ (
  .A(_0049_),
  .B1(_0622_),
  .B2(_0050_),
  .ZN(_0051_)
);

INV_X1 _1774_ (
  .A(_0051_),
  .ZN(_0052_)
);

OAI21_X1 _1775_ (
  .A(_0052_),
  .B1(_0619_),
  .B2(_0050_),
  .ZN(_0053_)
);

BUF_X2 _1776_ (
  .A(_1103_),
  .Z(_0054_)
);

XNOR2_X1 _1777_ (
  .A(_0053_),
  .B(_0054_),
  .ZN(_0055_)
);

NAND2_X1 _1778_ (
  .A1(_0055_),
  .A2(_0604_),
  .ZN(_0056_)
);

NAND2_X1 _1779_ (
  .A1(_0384_),
  .A2(_0581_),
  .ZN(_0057_)
);

NAND3_X1 _1780_ (
  .A1(_0056_),
  .A2(_0374_),
  .A3(_0057_),
  .ZN(_0058_)
);

INV_X1 _1781_ (
  .A(result[7]),
  .ZN(_0059_)
);

OAI21_X1 _1782_ (
  .A(_0058_),
  .B1(_0403_),
  .B2(_0059_),
  .ZN(_0026_)
);

NAND2_X1 _1783_ (
  .A1(_0385_),
  .A2(result[8]),
  .ZN(_0060_)
);

INV_X1 _1784_ (
  .A(_1102_),
  .ZN(_0061_)
);

INV_X1 _1785_ (
  .A(_0054_),
  .ZN(_0062_)
);

OAI21_X1 _1786_ (
  .A(_0061_),
  .B1(_0062_),
  .B2(_0047_),
  .ZN(_0063_)
);

INV_X1 _1787_ (
  .A(_0063_),
  .ZN(_0064_)
);

NAND2_X1 _1788_ (
  .A1(_0636_),
  .A2(_0054_),
  .ZN(_0065_)
);

OAI21_X1 _1789_ (
  .A(_0064_),
  .B1(_0632_),
  .B2(_0065_),
  .ZN(_0066_)
);

INV_X1 _1790_ (
  .A(_0066_),
  .ZN(_0067_)
);

NOR2_X1 _1791_ (
  .A1(_0634_),
  .A2(_0065_),
  .ZN(_0068_)
);

INV_X1 _1792_ (
  .A(_0068_),
  .ZN(_0069_)
);

OAI21_X1 _1793_ (
  .A(_0067_),
  .B1(_0633_),
  .B2(_0069_),
  .ZN(_0070_)
);

INV_X1 _1794_ (
  .A(_1105_),
  .ZN(_0071_)
);

XNOR2_X1 _1795_ (
  .A(_0070_),
  .B(_0071_),
  .ZN(_0072_)
);

OAI21_X1 _1796_ (
  .A(_0368_),
  .B1(_0072_),
  .B2(_0581_),
  .ZN(_0073_)
);

NOR2_X1 _1797_ (
  .A1(_0584_),
  .A2(\ext_mult_res[8] ),
  .ZN(_0074_)
);

OAI21_X1 _1798_ (
  .A(_0060_),
  .B1(_0073_),
  .B2(_0074_),
  .ZN(_0027_)
);

OAI21_X1 _1799_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[9] ),
  .ZN(_0075_)
);

INV_X1 _1800_ (
  .A(_0075_),
  .ZN(_0076_)
);

NAND2_X2 _1801_ (
  .A1(_0054_),
  .A2(_1105_),
  .ZN(_0077_)
);

INV_X1 _1802_ (
  .A(_0077_),
  .ZN(_0078_)
);

NAND2_X1 _1803_ (
  .A1(_0053_),
  .A2(_0078_),
  .ZN(_0079_)
);

INV_X1 _1804_ (
  .A(_1104_),
  .ZN(_0080_)
);

OAI21_X1 _1805_ (
  .A(_0080_),
  .B1(_0071_),
  .B2(_0061_),
  .ZN(_0081_)
);

INV_X1 _1806_ (
  .A(_0081_),
  .ZN(_0082_)
);

NAND2_X1 _1807_ (
  .A1(_0079_),
  .A2(_0082_),
  .ZN(_0083_)
);

INV_X1 _1808_ (
  .A(_1107_),
  .ZN(_0084_)
);

XNOR2_X1 _1809_ (
  .A(_0083_),
  .B(_0084_),
  .ZN(_0085_)
);

OAI21_X1 _1810_ (
  .A(_0076_),
  .B1(_0085_),
  .B2(_0581_),
  .ZN(_0086_)
);

NAND2_X1 _1811_ (
  .A1(_0387_),
  .A2(result[9]),
  .ZN(_0087_)
);

NAND2_X1 _1812_ (
  .A1(_0086_),
  .A2(_0087_),
  .ZN(_0028_)
);

NAND2_X1 _1813_ (
  .A1(_0385_),
  .A2(result[10]),
  .ZN(_0088_)
);

OAI21_X1 _1814_ (
  .A(_0632_),
  .B1(_0611_),
  .B2(_0634_),
  .ZN(_0089_)
);

NAND2_X1 _1815_ (
  .A1(_1105_),
  .A2(_1107_),
  .ZN(_0090_)
);

NOR2_X1 _1816_ (
  .A1(_0065_),
  .A2(_0090_),
  .ZN(_0091_)
);

NAND2_X1 _1817_ (
  .A1(_0089_),
  .A2(_0091_),
  .ZN(_0092_)
);

INV_X1 _1818_ (
  .A(_1106_),
  .ZN(_0093_)
);

OAI21_X1 _1819_ (
  .A(_0093_),
  .B1(_0084_),
  .B2(_0080_),
  .ZN(_0094_)
);

INV_X1 _1820_ (
  .A(_0094_),
  .ZN(_0095_)
);

OAI21_X1 _1821_ (
  .A(_0095_),
  .B1(_0064_),
  .B2(_0090_),
  .ZN(_0096_)
);

INV_X1 _1822_ (
  .A(_0096_),
  .ZN(_0097_)
);

NOR3_X1 _1823_ (
  .A1(_0634_),
  .A2(_0589_),
  .A3(_0609_),
  .ZN(_0098_)
);

INV_X1 _1824_ (
  .A(_0679_),
  .ZN(_0099_)
);

NAND3_X1 _1825_ (
  .A1(_0098_),
  .A2(_0099_),
  .A3(_0091_),
  .ZN(_0100_)
);

NAND3_X1 _1826_ (
  .A1(_0092_),
  .A2(_0097_),
  .A3(_0100_),
  .ZN(_0101_)
);

INV_X1 _1827_ (
  .A(_1109_),
  .ZN(_0102_)
);

XNOR2_X1 _1828_ (
  .A(_0101_),
  .B(_0102_),
  .ZN(_0103_)
);

NOR2_X1 _1829_ (
  .A1(_0103_),
  .A2(_0581_),
  .ZN(_0104_)
);

OAI21_X1 _1830_ (
  .A(_0368_),
  .B1(_0584_),
  .B2(\ext_mult_res[10] ),
  .ZN(_0105_)
);

OAI21_X1 _1831_ (
  .A(_0088_),
  .B1(_0104_),
  .B2(_0105_),
  .ZN(_0029_)
);

NAND2_X1 _1832_ (
  .A1(_0385_),
  .A2(result[11]),
  .ZN(_0106_)
);

NAND2_X1 _1833_ (
  .A1(_1107_),
  .A2(_1109_),
  .ZN(_0107_)
);

NOR2_X2 _1834_ (
  .A1(_0077_),
  .A2(_0107_),
  .ZN(_0108_)
);

NAND2_X1 _1835_ (
  .A1(_0051_),
  .A2(_0108_),
  .ZN(_0109_)
);

INV_X1 _1836_ (
  .A(_1108_),
  .ZN(_0110_)
);

OAI21_X1 _1837_ (
  .A(_0110_),
  .B1(_0102_),
  .B2(_0093_),
  .ZN(_0111_)
);

INV_X1 _1838_ (
  .A(_0111_),
  .ZN(_0112_)
);

OAI21_X1 _1839_ (
  .A(_0112_),
  .B1(_0082_),
  .B2(_0107_),
  .ZN(_0113_)
);

INV_X1 _1840_ (
  .A(_0113_),
  .ZN(_0114_)
);

NAND2_X1 _1841_ (
  .A1(_0109_),
  .A2(_0114_),
  .ZN(_0115_)
);

INV_X1 _1842_ (
  .A(_0115_),
  .ZN(_0116_)
);

NAND4_X1 _1843_ (
  .A1(_0108_),
  .A2(_0618_),
  .A3(_0636_),
  .A4(_0624_),
  .ZN(_0117_)
);

INV_X1 _1844_ (
  .A(_0117_),
  .ZN(_0118_)
);

INV_X1 _1845_ (
  .A(_0602_),
  .ZN(_0119_)
);

NAND2_X1 _1846_ (
  .A1(_0118_),
  .A2(_0119_),
  .ZN(_0120_)
);

NAND2_X1 _1847_ (
  .A1(_0116_),
  .A2(_0120_),
  .ZN(_0121_)
);

INV_X1 _1848_ (
  .A(_1111_),
  .ZN(_0122_)
);

NAND2_X1 _1849_ (
  .A1(_0121_),
  .A2(_0122_),
  .ZN(_0123_)
);

NAND3_X1 _1850_ (
  .A1(_0116_),
  .A2(_1111_),
  .A3(_0120_),
  .ZN(_0124_)
);

NAND3_X1 _1851_ (
  .A1(_0123_),
  .A2(_0124_),
  .A3(_0604_),
  .ZN(_0125_)
);

NAND2_X1 _1852_ (
  .A1(_0125_),
  .A2(_0374_),
  .ZN(_0126_)
);

NOR2_X1 _1853_ (
  .A1(_0584_),
  .A2(\ext_mult_res[11] ),
  .ZN(_0127_)
);

OAI21_X1 _1854_ (
  .A(_0106_),
  .B1(_0126_),
  .B2(_0127_),
  .ZN(_0030_)
);

NAND2_X1 _1855_ (
  .A1(_0385_),
  .A2(result[12]),
  .ZN(_0128_)
);

NAND2_X1 _1856_ (
  .A1(_1109_),
  .A2(_1111_),
  .ZN(_0129_)
);

NOR2_X1 _1857_ (
  .A1(_0090_),
  .A2(_0129_),
  .ZN(_0130_)
);

NAND2_X1 _1858_ (
  .A1(_0066_),
  .A2(_0130_),
  .ZN(_0131_)
);

INV_X1 _1859_ (
  .A(_1110_),
  .ZN(_0132_)
);

OAI21_X1 _1860_ (
  .A(_0132_),
  .B1(_0122_),
  .B2(_0110_),
  .ZN(_0133_)
);

INV_X1 _1861_ (
  .A(_0133_),
  .ZN(_0134_)
);

OAI21_X1 _1862_ (
  .A(_0134_),
  .B1(_0095_),
  .B2(_0129_),
  .ZN(_0135_)
);

INV_X1 _1863_ (
  .A(_0135_),
  .ZN(_0136_)
);

NAND2_X1 _1864_ (
  .A1(_0131_),
  .A2(_0136_),
  .ZN(_0137_)
);

INV_X1 _1865_ (
  .A(_0137_),
  .ZN(_0138_)
);

NAND2_X1 _1866_ (
  .A1(_0068_),
  .A2(_0130_),
  .ZN(_0139_)
);

INV_X1 _1867_ (
  .A(_0139_),
  .ZN(_0140_)
);

NAND2_X1 _1868_ (
  .A1(_0612_),
  .A2(_0140_),
  .ZN(_0141_)
);

NAND2_X1 _1869_ (
  .A1(_0138_),
  .A2(_0141_),
  .ZN(_0142_)
);

INV_X1 _1870_ (
  .A(_1113_),
  .ZN(_0143_)
);

NAND2_X1 _1871_ (
  .A1(_0142_),
  .A2(_0143_),
  .ZN(_0144_)
);

NAND3_X1 _1872_ (
  .A1(_0138_),
  .A2(_1113_),
  .A3(_0141_),
  .ZN(_0145_)
);

AND3_X1 _1873_ (
  .A1(_0144_),
  .A2(_0145_),
  .A3(_0594_),
  .ZN(_0146_)
);

OAI21_X1 _1874_ (
  .A(_0368_),
  .B1(_0584_),
  .B2(\ext_mult_res[12] ),
  .ZN(_0147_)
);

OAI21_X1 _1875_ (
  .A(_0128_),
  .B1(_0146_),
  .B2(_0147_),
  .ZN(_0031_)
);

NAND2_X1 _1876_ (
  .A1(_0385_),
  .A2(result[13]),
  .ZN(_0148_)
);

NAND2_X1 _1877_ (
  .A1(_0048_),
  .A2(_0078_),
  .ZN(_0149_)
);

NAND2_X1 _1878_ (
  .A1(_0082_),
  .A2(_0149_),
  .ZN(_0150_)
);

NAND2_X1 _1879_ (
  .A1(_1111_),
  .A2(_1113_),
  .ZN(_0151_)
);

NOR2_X1 _1880_ (
  .A1(_0107_),
  .A2(_0151_),
  .ZN(_0152_)
);

NAND2_X1 _1881_ (
  .A1(_0150_),
  .A2(_0152_),
  .ZN(_0153_)
);

INV_X1 _1882_ (
  .A(_0151_),
  .ZN(_0154_)
);

NAND2_X1 _1883_ (
  .A1(_0111_),
  .A2(_0154_),
  .ZN(_0155_)
);

INV_X1 _1884_ (
  .A(_1112_),
  .ZN(_0156_)
);

OAI21_X1 _1885_ (
  .A(_0156_),
  .B1(_0143_),
  .B2(_0132_),
  .ZN(_0157_)
);

INV_X1 _1886_ (
  .A(_0157_),
  .ZN(_0158_)
);

NAND2_X1 _1887_ (
  .A1(_0155_),
  .A2(_0158_),
  .ZN(_0159_)
);

INV_X1 _1888_ (
  .A(_0159_),
  .ZN(_0160_)
);

NAND2_X1 _1889_ (
  .A1(_0153_),
  .A2(_0160_),
  .ZN(_0161_)
);

INV_X1 _1890_ (
  .A(_0161_),
  .ZN(_0162_)
);

INV_X1 _1891_ (
  .A(_0623_),
  .ZN(_0163_)
);

NOR2_X2 _1892_ (
  .A1(_0050_),
  .A2(_0077_),
  .ZN(_0164_)
);

NAND2_X1 _1893_ (
  .A1(_0164_),
  .A2(_0152_),
  .ZN(_0165_)
);

OAI21_X1 _1894_ (
  .A(_0162_),
  .B1(_0163_),
  .B2(_0165_),
  .ZN(_0166_)
);

INV_X1 _1895_ (
  .A(_1115_),
  .ZN(_0167_)
);

XNOR2_X1 _1896_ (
  .A(_0166_),
  .B(_0167_),
  .ZN(_0168_)
);

NOR2_X1 _1897_ (
  .A1(_0168_),
  .A2(_0581_),
  .ZN(_0169_)
);

OAI21_X1 _1898_ (
  .A(_0368_),
  .B1(_0604_),
  .B2(\ext_mult_res[13] ),
  .ZN(_0170_)
);

OAI21_X1 _1899_ (
  .A(_0148_),
  .B1(_0169_),
  .B2(_0170_),
  .ZN(_0032_)
);

NAND2_X1 _1900_ (
  .A1(_1113_),
  .A2(_1115_),
  .ZN(_0171_)
);

NOR2_X1 _1901_ (
  .A1(_0129_),
  .A2(_0171_),
  .ZN(_0172_)
);

NAND3_X1 _1902_ (
  .A1(_0635_),
  .A2(_0091_),
  .A3(_0172_),
  .ZN(_0173_)
);

INV_X1 _1903_ (
  .A(_1114_),
  .ZN(_0174_)
);

OAI21_X1 _1904_ (
  .A(_0174_),
  .B1(_0167_),
  .B2(_0156_),
  .ZN(_0175_)
);

INV_X1 _1905_ (
  .A(_0175_),
  .ZN(_0176_)
);

OAI21_X1 _1906_ (
  .A(_0176_),
  .B1(_0134_),
  .B2(_0171_),
  .ZN(_0177_)
);

AOI21_X1 _1907_ (
  .A(_0177_),
  .B1(_0172_),
  .B2(_0096_),
  .ZN(_0178_)
);

NAND2_X1 _1908_ (
  .A1(_0173_),
  .A2(_0178_),
  .ZN(_0179_)
);

INV_X1 _1909_ (
  .A(_1117_),
  .ZN(_0180_)
);

NAND2_X1 _1910_ (
  .A1(_0179_),
  .A2(_0180_),
  .ZN(_0181_)
);

NAND3_X1 _1911_ (
  .A1(_0173_),
  .A2(_1117_),
  .A3(_0178_),
  .ZN(_0182_)
);

NAND3_X1 _1912_ (
  .A1(_0181_),
  .A2(_0182_),
  .A3(_0604_),
  .ZN(_0183_)
);

OAI21_X1 _1913_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[14] ),
  .ZN(_0184_)
);

INV_X1 _1914_ (
  .A(_0184_),
  .ZN(_0185_)
);

NAND2_X1 _1915_ (
  .A1(_0183_),
  .A2(_0185_),
  .ZN(_0186_)
);

NAND2_X1 _1916_ (
  .A1(_0387_),
  .A2(result[14]),
  .ZN(_0187_)
);

NAND2_X1 _1917_ (
  .A1(_0186_),
  .A2(_0187_),
  .ZN(_0033_)
);

NAND2_X1 _1918_ (
  .A1(_1115_),
  .A2(_1117_),
  .ZN(_0188_)
);

NOR2_X1 _1919_ (
  .A1(_0151_),
  .A2(_0188_),
  .ZN(_0189_)
);

NAND3_X1 _1920_ (
  .A1(_0053_),
  .A2(_0108_),
  .A3(_0189_),
  .ZN(_0190_)
);

INV_X1 _1921_ (
  .A(_1116_),
  .ZN(_0191_)
);

OAI21_X1 _1922_ (
  .A(_0191_),
  .B1(_0180_),
  .B2(_0174_),
  .ZN(_0192_)
);

INV_X1 _1923_ (
  .A(_0192_),
  .ZN(_0193_)
);

OAI21_X1 _1924_ (
  .A(_0193_),
  .B1(_0158_),
  .B2(_0188_),
  .ZN(_0194_)
);

AOI21_X1 _1925_ (
  .A(_0194_),
  .B1(_0189_),
  .B2(_0113_),
  .ZN(_0195_)
);

NAND2_X1 _1926_ (
  .A1(_0190_),
  .A2(_0195_),
  .ZN(_0196_)
);

INV_X1 _1927_ (
  .A(_1119_),
  .ZN(_0197_)
);

NAND2_X1 _1928_ (
  .A1(_0196_),
  .A2(_0197_),
  .ZN(_0198_)
);

NAND3_X1 _1929_ (
  .A1(_0190_),
  .A2(_1119_),
  .A3(_0195_),
  .ZN(_0199_)
);

NAND3_X1 _1930_ (
  .A1(_0198_),
  .A2(_0199_),
  .A3(_0604_),
  .ZN(_0200_)
);

OAI21_X1 _1931_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[15] ),
  .ZN(_0201_)
);

INV_X1 _1932_ (
  .A(_0201_),
  .ZN(_0202_)
);

NAND2_X1 _1933_ (
  .A1(_0200_),
  .A2(_0202_),
  .ZN(_0203_)
);

NAND2_X1 _1934_ (
  .A1(_0387_),
  .A2(result[15]),
  .ZN(_0204_)
);

NAND2_X1 _1935_ (
  .A1(_0203_),
  .A2(_0204_),
  .ZN(_0034_)
);

OAI21_X1 _1936_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[16] ),
  .ZN(_0205_)
);

INV_X1 _1937_ (
  .A(_0205_),
  .ZN(_0206_)
);

NAND2_X1 _1938_ (
  .A1(_1117_),
  .A2(_1119_),
  .ZN(_0207_)
);

NOR2_X1 _1939_ (
  .A1(_0171_),
  .A2(_0207_),
  .ZN(_0208_)
);

NAND3_X1 _1940_ (
  .A1(_0070_),
  .A2(_0130_),
  .A3(_0208_),
  .ZN(_0209_)
);

BUF_X2 _1941_ (
  .A(_1121_),
  .Z(_0210_)
);

INV_X1 _1942_ (
  .A(_1118_),
  .ZN(_0211_)
);

OAI21_X1 _1943_ (
  .A(_0211_),
  .B1(_0197_),
  .B2(_0191_),
  .ZN(_0212_)
);

INV_X1 _1944_ (
  .A(_0212_),
  .ZN(_0213_)
);

OAI21_X1 _1945_ (
  .A(_0213_),
  .B1(_0176_),
  .B2(_0207_),
  .ZN(_0214_)
);

AOI21_X1 _1946_ (
  .A(_0214_),
  .B1(_0208_),
  .B2(_0135_),
  .ZN(_0215_)
);

NAND3_X1 _1947_ (
  .A1(_0209_),
  .A2(_0210_),
  .A3(_0215_),
  .ZN(_0216_)
);

NAND2_X1 _1948_ (
  .A1(_0216_),
  .A2(_0604_),
  .ZN(_0217_)
);

AOI21_X1 _1949_ (
  .A(_0210_),
  .B1(_0209_),
  .B2(_0215_),
  .ZN(_0218_)
);

OAI21_X1 _1950_ (
  .A(_0206_),
  .B1(_0217_),
  .B2(_0218_),
  .ZN(_0219_)
);

NAND2_X1 _1951_ (
  .A1(_0387_),
  .A2(result[16]),
  .ZN(_0220_)
);

NAND2_X1 _1952_ (
  .A1(_0219_),
  .A2(_0220_),
  .ZN(_0035_)
);

OAI21_X1 _1953_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[17] ),
  .ZN(_0221_)
);

INV_X1 _1954_ (
  .A(_0221_),
  .ZN(_0222_)
);

OAI21_X1 _1955_ (
  .A(_0599_),
  .B1(_0589_),
  .B2(_0598_),
  .ZN(_0223_)
);

INV_X1 _1956_ (
  .A(_0223_),
  .ZN(_0224_)
);

OAI21_X1 _1957_ (
  .A(_0622_),
  .B1(_0224_),
  .B2(_0617_),
  .ZN(_0225_)
);

NAND2_X1 _1958_ (
  .A1(_0225_),
  .A2(_0164_),
  .ZN(_0226_)
);

INV_X1 _1959_ (
  .A(_0150_),
  .ZN(_0227_)
);

NAND2_X1 _1960_ (
  .A1(_0226_),
  .A2(_0227_),
  .ZN(_0228_)
);

NAND2_X2 _1961_ (
  .A1(_1119_),
  .A2(_0210_),
  .ZN(_0229_)
);

NOR2_X2 _1962_ (
  .A1(_0188_),
  .A2(_0229_),
  .ZN(_0230_)
);

AND2_X1 _1963_ (
  .A1(_0152_),
  .A2(_0230_),
  .ZN(_0231_)
);

NAND2_X1 _1964_ (
  .A1(_0228_),
  .A2(_0231_),
  .ZN(_0232_)
);

INV_X1 _1965_ (
  .A(_0229_),
  .ZN(_0233_)
);

NAND2_X1 _1966_ (
  .A1(_0192_),
  .A2(_0233_),
  .ZN(_0234_)
);

INV_X1 _1967_ (
  .A(_1120_),
  .ZN(_0235_)
);

INV_X1 _1968_ (
  .A(_0210_),
  .ZN(_0236_)
);

OAI21_X1 _1969_ (
  .A(_0235_),
  .B1(_0236_),
  .B2(_0211_),
  .ZN(_0237_)
);

INV_X1 _1970_ (
  .A(_0237_),
  .ZN(_0238_)
);

NAND2_X1 _1971_ (
  .A1(_0234_),
  .A2(_0238_),
  .ZN(_0239_)
);

AOI21_X1 _1972_ (
  .A(_0239_),
  .B1(_0230_),
  .B2(_0159_),
  .ZN(_0240_)
);

AND3_X1 _1973_ (
  .A1(_0618_),
  .A2(_1091_),
  .A3(_1093_),
  .ZN(_0241_)
);

NAND4_X1 _1974_ (
  .A1(_0231_),
  .A2(_0241_),
  .A3(_0164_),
  .A4(_1088_),
  .ZN(_0242_)
);

NAND3_X1 _1975_ (
  .A1(_0232_),
  .A2(_0240_),
  .A3(_0242_),
  .ZN(_0243_)
);

INV_X1 _1976_ (
  .A(_1123_),
  .ZN(_0244_)
);

NAND2_X1 _1977_ (
  .A1(_0243_),
  .A2(_0244_),
  .ZN(_0245_)
);

NAND2_X1 _1978_ (
  .A1(_0245_),
  .A2(_0604_),
  .ZN(_0246_)
);

NOR2_X1 _1979_ (
  .A1(_0243_),
  .A2(_0244_),
  .ZN(_0247_)
);

OAI21_X1 _1980_ (
  .A(_0222_),
  .B1(_0246_),
  .B2(_0247_),
  .ZN(_0248_)
);

NAND2_X1 _1981_ (
  .A1(_0387_),
  .A2(result[17]),
  .ZN(_0249_)
);

NAND2_X1 _1982_ (
  .A1(_0248_),
  .A2(_0249_),
  .ZN(_0036_)
);

NOR2_X1 _1983_ (
  .A1(_0368_),
  .A2(result[18]),
  .ZN(_0250_)
);

NAND2_X1 _1984_ (
  .A1(_0092_),
  .A2(_0097_),
  .ZN(_0251_)
);

NAND2_X1 _1985_ (
  .A1(_0210_),
  .A2(_1123_),
  .ZN(_0252_)
);

NOR2_X1 _1986_ (
  .A1(_0207_),
  .A2(_0252_),
  .ZN(_0253_)
);

AND2_X1 _1987_ (
  .A1(_0172_),
  .A2(_0253_),
  .ZN(_0254_)
);

NAND2_X1 _1988_ (
  .A1(_0251_),
  .A2(_0254_),
  .ZN(_0255_)
);

INV_X1 _1989_ (
  .A(_1122_),
  .ZN(_0256_)
);

OAI21_X1 _1990_ (
  .A(_0256_),
  .B1(_0244_),
  .B2(_0235_),
  .ZN(_0257_)
);

INV_X1 _1991_ (
  .A(_0257_),
  .ZN(_0258_)
);

OAI21_X1 _1992_ (
  .A(_0258_),
  .B1(_0213_),
  .B2(_0252_),
  .ZN(_0259_)
);

AOI21_X1 _1993_ (
  .A(_0259_),
  .B1(_0253_),
  .B2(_0177_),
  .ZN(_0260_)
);

NAND4_X1 _1994_ (
  .A1(_0254_),
  .A2(_0091_),
  .A3(_0098_),
  .A4(_0099_),
  .ZN(_0261_)
);

NAND3_X1 _1995_ (
  .A1(_0255_),
  .A2(_0260_),
  .A3(_0261_),
  .ZN(_0262_)
);

NAND2_X1 _1996_ (
  .A1(_0262_),
  .A2(_1125_),
  .ZN(_0263_)
);

INV_X1 _1997_ (
  .A(_1125_),
  .ZN(_0264_)
);

NAND4_X1 _1998_ (
  .A1(_0255_),
  .A2(_0260_),
  .A3(_0264_),
  .A4(_0261_),
  .ZN(_0265_)
);

NAND3_X1 _1999_ (
  .A1(_0263_),
  .A2(_0265_),
  .A3(_0584_),
  .ZN(_0266_)
);

NAND2_X1 _2000_ (
  .A1(_0581_),
  .A2(\ext_mult_res[18] ),
  .ZN(_0267_)
);

NAND2_X1 _2001_ (
  .A1(_0267_),
  .A2(_0371_),
  .ZN(_0268_)
);

INV_X1 _2002_ (
  .A(_0268_),
  .ZN(_0269_)
);

AOI21_X1 _2003_ (
  .A(_0250_),
  .B1(_0266_),
  .B2(_0269_),
  .ZN(_0037_)
);

NOR2_X1 _2004_ (
  .A1(_0368_),
  .A2(result[19]),
  .ZN(_0270_)
);

NAND2_X1 _2005_ (
  .A1(_1123_),
  .A2(_1125_),
  .ZN(_0271_)
);

NOR2_X1 _2006_ (
  .A1(_0229_),
  .A2(_0271_),
  .ZN(_0272_)
);

AND2_X1 _2007_ (
  .A1(_0189_),
  .A2(_0272_),
  .ZN(_0273_)
);

NAND2_X1 _2008_ (
  .A1(_0115_),
  .A2(_0273_),
  .ZN(_0274_)
);

INV_X1 _2009_ (
  .A(_1124_),
  .ZN(_0275_)
);

OAI21_X1 _2010_ (
  .A(_0275_),
  .B1(_0264_),
  .B2(_0256_),
  .ZN(_0276_)
);

INV_X1 _2011_ (
  .A(_0276_),
  .ZN(_0277_)
);

OAI21_X1 _2012_ (
  .A(_0277_),
  .B1(_0238_),
  .B2(_0271_),
  .ZN(_0278_)
);

AOI21_X1 _2013_ (
  .A(_0278_),
  .B1(_0272_),
  .B2(_0194_),
  .ZN(_0279_)
);

NAND3_X1 _2014_ (
  .A1(_0118_),
  .A2(_0119_),
  .A3(_0273_),
  .ZN(_0280_)
);

NAND3_X1 _2015_ (
  .A1(_0274_),
  .A2(_0279_),
  .A3(_0280_),
  .ZN(_0281_)
);

NAND2_X1 _2016_ (
  .A1(_0281_),
  .A2(_1127_),
  .ZN(_0282_)
);

INV_X1 _2017_ (
  .A(_1127_),
  .ZN(_0283_)
);

NAND4_X1 _2018_ (
  .A1(_0274_),
  .A2(_0279_),
  .A3(_0283_),
  .A4(_0280_),
  .ZN(_0284_)
);

NAND3_X1 _2019_ (
  .A1(_0282_),
  .A2(_0284_),
  .A3(_0584_),
  .ZN(_0285_)
);

AOI21_X1 _2020_ (
  .A(_0270_),
  .B1(_0285_),
  .B2(_0269_),
  .ZN(_0038_)
);

NOR2_X1 _2021_ (
  .A1(_0368_),
  .A2(result[20]),
  .ZN(_0286_)
);

NAND2_X1 _2022_ (
  .A1(_1125_),
  .A2(_1127_),
  .ZN(_0287_)
);

NOR2_X1 _2023_ (
  .A1(_0252_),
  .A2(_0287_),
  .ZN(_0288_)
);

AND2_X1 _2024_ (
  .A1(_0208_),
  .A2(_0288_),
  .ZN(_0289_)
);

NAND2_X1 _2025_ (
  .A1(_0137_),
  .A2(_0289_),
  .ZN(_0290_)
);

INV_X1 _2026_ (
  .A(_1126_),
  .ZN(_0291_)
);

OAI21_X1 _2027_ (
  .A(_0291_),
  .B1(_0283_),
  .B2(_0275_),
  .ZN(_0292_)
);

INV_X1 _2028_ (
  .A(_0292_),
  .ZN(_0293_)
);

OAI21_X1 _2029_ (
  .A(_0293_),
  .B1(_0258_),
  .B2(_0287_),
  .ZN(_0294_)
);

AOI21_X1 _2030_ (
  .A(_0294_),
  .B1(_0288_),
  .B2(_0214_),
  .ZN(_0295_)
);

NAND3_X1 _2031_ (
  .A1(_0612_),
  .A2(_0140_),
  .A3(_0289_),
  .ZN(_0296_)
);

NAND3_X1 _2032_ (
  .A1(_0290_),
  .A2(_0295_),
  .A3(_0296_),
  .ZN(_0297_)
);

NAND2_X1 _2033_ (
  .A1(_0297_),
  .A2(_1129_),
  .ZN(_0298_)
);

INV_X1 _2034_ (
  .A(_1129_),
  .ZN(_0299_)
);

NAND4_X1 _2035_ (
  .A1(_0290_),
  .A2(_0295_),
  .A3(_0299_),
  .A4(_0296_),
  .ZN(_0300_)
);

NAND3_X1 _2036_ (
  .A1(_0298_),
  .A2(_0300_),
  .A3(_0584_),
  .ZN(_0301_)
);

AOI21_X1 _2037_ (
  .A(_0286_),
  .B1(_0301_),
  .B2(_0269_),
  .ZN(_0039_)
);

NAND2_X1 _2038_ (
  .A1(_1127_),
  .A2(_1129_),
  .ZN(_0302_)
);

NOR2_X1 _2039_ (
  .A1(_0271_),
  .A2(_0302_),
  .ZN(_0303_)
);

NAND2_X1 _2040_ (
  .A1(_0230_),
  .A2(_0303_),
  .ZN(_0304_)
);

INV_X1 _2041_ (
  .A(_0304_),
  .ZN(_0305_)
);

NAND2_X1 _2042_ (
  .A1(_0161_),
  .A2(_0305_),
  .ZN(_0306_)
);

INV_X1 _2043_ (
  .A(_0303_),
  .ZN(_0307_)
);

AOI21_X1 _2044_ (
  .A(_0307_),
  .B1(_0234_),
  .B2(_0238_),
  .ZN(_0308_)
);

INV_X1 _2045_ (
  .A(_1128_),
  .ZN(_0309_)
);

OAI21_X1 _2046_ (
  .A(_0309_),
  .B1(_0299_),
  .B2(_0291_),
  .ZN(_0310_)
);

INV_X1 _2047_ (
  .A(_0310_),
  .ZN(_0311_)
);

OAI21_X1 _2048_ (
  .A(_0311_),
  .B1(_0277_),
  .B2(_0302_),
  .ZN(_0312_)
);

NOR2_X1 _2049_ (
  .A1(_0308_),
  .A2(_0312_),
  .ZN(_0313_)
);

NOR2_X1 _2050_ (
  .A1(_0165_),
  .A2(_0304_),
  .ZN(_0314_)
);

NAND2_X1 _2051_ (
  .A1(_0623_),
  .A2(_0314_),
  .ZN(_0315_)
);

XOR2_X1 _2052_ (
  .A(\ext_mult_res[18] ),
  .B(result[21]),
  .Z(_0316_)
);

NAND4_X1 _2053_ (
  .A1(_0306_),
  .A2(_0313_),
  .A3(_0315_),
  .A4(_0316_),
  .ZN(_0317_)
);

NAND3_X1 _2054_ (
  .A1(_0306_),
  .A2(_0313_),
  .A3(_0315_),
  .ZN(_0318_)
);

INV_X1 _2055_ (
  .A(_0316_),
  .ZN(_0319_)
);

NAND2_X1 _2056_ (
  .A1(_0318_),
  .A2(_0319_),
  .ZN(_0320_)
);

NAND2_X1 _2057_ (
  .A1(_0317_),
  .A2(_0320_),
  .ZN(_0321_)
);

NAND2_X1 _2058_ (
  .A1(_0321_),
  .A2(_0594_),
  .ZN(_0322_)
);

NAND2_X1 _2059_ (
  .A1(_0322_),
  .A2(_0267_),
  .ZN(_0323_)
);

NAND2_X1 _2060_ (
  .A1(_0323_),
  .A2(_0372_),
  .ZN(_0324_)
);

NAND2_X1 _2061_ (
  .A1(_0387_),
  .A2(result[21]),
  .ZN(_0325_)
);

NAND2_X1 _2062_ (
  .A1(_0324_),
  .A2(_0325_),
  .ZN(_0040_)
);

FA_X1 _2063_ (
  .A(_0676_),
  .B(_0677_),
  .CI(_0678_),
  .CO(_0679_),
  .S(_0680_)
);

FA_X1 _2064_ (
  .A(_0681_),
  .B(_0682_),
  .CI(_0683_),
  .CO(_0684_),
  .S(_0685_)
);

FA_X1 _2065_ (
  .A(_0686_),
  .B(_0687_),
  .CI(_0688_),
  .CO(_0689_),
  .S(_0690_)
);

FA_X1 _2066_ (
  .A(_0690_),
  .B(_0684_),
  .CI(_0691_),
  .CO(_0692_),
  .S(_0693_)
);

FA_X1 _2067_ (
  .A(_0694_),
  .B(_0695_),
  .CI(_0696_),
  .CO(_0697_),
  .S(_0698_)
);

FA_X1 _2068_ (
  .A(_0698_),
  .B(_0699_),
  .CI(_0700_),
  .CO(_0701_),
  .S(_0702_)
);

FA_X1 _2069_ (
  .A(_0703_),
  .B(_0704_),
  .CI(_0705_),
  .CO(_0706_),
  .S(_0707_)
);

FA_X1 _2070_ (
  .A(_0708_),
  .B(_0709_),
  .CI(_0710_),
  .CO(_0711_),
  .S(_0712_)
);

FA_X1 _2071_ (
  .A(_0707_),
  .B(_0697_),
  .CI(_0712_),
  .CO(_0713_),
  .S(_0714_)
);

FA_X1 _2072_ (
  .A(_0715_),
  .B(_0716_),
  .CI(_0717_),
  .CO(_0718_),
  .S(_0719_)
);

FA_X1 _2073_ (
  .A(_0720_),
  .B(_0721_),
  .CI(_0722_),
  .CO(_0723_),
  .S(_0724_)
);

FA_X1 _2074_ (
  .A(_0725_),
  .B(_0726_),
  .CI(_0727_),
  .CO(_0728_),
  .S(_0729_)
);

FA_X1 _2075_ (
  .A(_0724_),
  .B(_0706_),
  .CI(_0729_),
  .CO(_0730_),
  .S(_0731_)
);

FA_X1 _2076_ (
  .A(_0731_),
  .B(_0713_),
  .CI(_0732_),
  .CO(_0733_),
  .S(_0734_)
);

FA_X1 _2077_ (
  .A(_0735_),
  .B(_0736_),
  .CI(_0737_),
  .CO(_0738_),
  .S(_0739_)
);

FA_X1 _2078_ (
  .A(_0740_),
  .B(_0741_),
  .CI(_0742_),
  .CO(_0743_),
  .S(_0744_)
);

FA_X1 _2079_ (
  .A(_0744_),
  .B(_0739_),
  .CI(_0745_),
  .CO(_0746_),
  .S(_0747_)
);

FA_X1 _2080_ (
  .A(_0748_),
  .B(_0749_),
  .CI(_0750_),
  .CO(_0751_),
  .S(_0752_)
);

FA_X1 _2081_ (
  .A(_0753_),
  .B(_0754_),
  .CI(_0755_),
  .CO(_0756_),
  .S(_0757_)
);

FA_X1 _2082_ (
  .A(_0758_),
  .B(_0759_),
  .CI(_0760_),
  .CO(_0761_),
  .S(_0762_)
);

FA_X1 _2083_ (
  .A(_0765_),
  .B(_0766_),
  .CI(_0767_),
  .CO(_0768_),
  .S(_0769_)
);

FA_X1 _2084_ (
  .A(_0770_),
  .B(_0747_),
  .CI(_0771_),
  .CO(_0772_),
  .S(_0773_)
);

FA_X1 _2085_ (
  .A(_0757_),
  .B(_0774_),
  .CI(_0775_),
  .CO(_0776_),
  .S(_0777_)
);

FA_X1 _2086_ (
  .A(_0778_),
  .B(_0779_),
  .CI(_0780_),
  .CO(_0781_),
  .S(_0782_)
);

FA_X1 _2087_ (
  .A(_0777_),
  .B(_0730_),
  .CI(_0784_),
  .CO(_0783_),
  .S(_0785_)
);

FA_X1 _2088_ (
  .A(_0786_),
  .B(_0733_),
  .CI(_0787_),
  .CO(_0788_),
  .S(_0789_)
);

FA_X1 _2089_ (
  .A(_0790_),
  .B(_0791_),
  .CI(_0792_),
  .CO(_0793_),
  .S(_0794_)
);

FA_X1 _2090_ (
  .A(_0795_),
  .B(_0796_),
  .CI(_0797_),
  .CO(_0798_),
  .S(_0799_)
);

FA_X1 _2091_ (
  .A(_0800_),
  .B(_0801_),
  .CI(_0802_),
  .CO(_0803_),
  .S(_0804_)
);

FA_X1 _2092_ (
  .A(_0799_),
  .B(_0738_),
  .CI(_0804_),
  .CO(_0805_),
  .S(_0806_)
);

FA_X1 _2093_ (
  .A(_0759_),
  .B(_0807_),
  .CI(_0808_),
  .CO(_0809_),
  .S(_0810_)
);

FA_X1 _2094_ (
  .A(_0811_),
  .B(_0812_),
  .CI(_0813_),
  .CO(_0814_),
  .S(_0815_)
);

FA_X1 _2095_ (
  .A(_0806_),
  .B(_0746_),
  .CI(_0815_),
  .CO(_0816_),
  .S(_0817_)
);

FA_X1 _2096_ (
  .A(_0817_),
  .B(_0772_),
  .CI(_0818_),
  .CO(_0819_),
  .S(_0820_)
);

FA_X1 _2097_ (
  .A(_0821_),
  .B(_0822_),
  .CI(_0823_),
  .CO(_0824_),
  .S(_0825_)
);

FA_X1 _2098_ (
  .A(_0826_),
  .B(_0827_),
  .CI(_0828_),
  .CO(_0829_),
  .S(_0830_)
);

FA_X1 _2099_ (
  .A(_0825_),
  .B(_0798_),
  .CI(_0830_),
  .CO(_0831_),
  .S(_0832_)
);

FA_X1 _2100_ (
  .A(_0833_),
  .B(_0834_),
  .CI(_0808_),
  .CO(_0835_),
  .S(_0836_)
);

FA_X1 _2101_ (
  .A(_0837_),
  .B(_0838_),
  .CI(_0839_),
  .CO(_0840_),
  .S(_0841_)
);

FA_X1 _2102_ (
  .A(_0841_),
  .B(_0832_),
  .CI(_0805_),
  .CO(_0842_),
  .S(_0843_)
);

FA_X1 _2103_ (
  .A(_0816_),
  .B(_0843_),
  .CI(_0844_),
  .CO(_0845_),
  .S(_0846_)
);

FA_X1 _2104_ (
  .A(_0847_),
  .B(_0848_),
  .CI(_0849_),
  .CO(_0850_),
  .S(_0851_)
);

FA_X1 _2105_ (
  .A(_0852_),
  .B(_0853_),
  .CI(_0854_),
  .CO(_0855_),
  .S(_0856_)
);

FA_X1 _2106_ (
  .A(_0857_),
  .B(_0858_),
  .CI(_0859_),
  .CO(_0860_),
  .S(_0861_)
);

FA_X1 _2107_ (
  .A(_0862_),
  .B(_0824_),
  .CI(_0861_),
  .CO(_0863_),
  .S(_0864_)
);

FA_X1 _2108_ (
  .A(_0833_),
  .B(_0865_),
  .CI(_0866_),
  .CO(_0867_),
  .S(_0868_)
);

FA_X1 _2109_ (
  .A(_0829_),
  .B(_0868_),
  .CI(_0835_),
  .CO(_0869_),
  .S(_0870_)
);

FA_X1 _2110_ (
  .A(_0864_),
  .B(_0831_),
  .CI(_0870_),
  .CO(_0871_),
  .S(_0872_)
);

FA_X1 _2111_ (
  .A(_0763_),
  .B(_0764_),
  .CI(_0873_),
  .CO(_0874_),
  .S(_0875_)
);

FA_X1 _2112_ (
  .A(_0872_),
  .B(_0842_),
  .CI(_0876_),
  .CO(_0877_),
  .S(_0878_)
);

FA_X1 _2113_ (
  .A(_0878_),
  .B(_0845_),
  .CI(_0879_),
  .CO(_0880_),
  .S(_0881_)
);

FA_X1 _2114_ (
  .A(_0852_),
  .B(_0882_),
  .CI(_0854_),
  .CO(_0883_),
  .S(_0884_)
);

FA_X1 _2115_ (
  .A(_0885_),
  .B(_0886_),
  .CI(_0887_),
  .CO(_0888_),
  .S(_0889_)
);

FA_X1 _2116_ (
  .A(_0890_),
  .B(_0891_),
  .CI(_0889_),
  .CO(_0892_),
  .S(_0893_)
);

FA_X1 _2117_ (
  .A(_0866_),
  .B(_0894_),
  .CI(_0895_),
  .CO(_0896_),
  .S(_0897_)
);

FA_X1 _2118_ (
  .A(_0860_),
  .B(_0897_),
  .CI(_0867_),
  .CO(_0898_),
  .S(_0899_)
);

FA_X1 _2119_ (
  .A(_0893_),
  .B(_0863_),
  .CI(_0899_),
  .CO(_0900_),
  .S(_0901_)
);

FA_X1 _2120_ (
  .A(_0759_),
  .B(_0833_),
  .CI(_0808_),
  .CO(_0902_),
  .S(_0903_)
);

FA_X1 _2121_ (
  .A(_0760_),
  .B(_0904_),
  .CI(_0905_),
  .CO(_0906_),
  .S(_0907_)
);

FA_X1 _2122_ (
  .A(_0908_),
  .B(_0909_),
  .CI(_0910_),
  .CO(_0911_),
  .S(_0912_)
);

FA_X1 _2123_ (
  .A(_0901_),
  .B(_0871_),
  .CI(_0913_),
  .CO(_0914_),
  .S(_0915_)
);

FA_X1 _2124_ (
  .A(_0915_),
  .B(_0877_),
  .CI(_0916_),
  .CO(_0917_),
  .S(_0918_)
);

FA_X1 _2125_ (
  .A(_0919_),
  .B(_0920_),
  .CI(_0921_),
  .CO(_0922_),
  .S(_0923_)
);

FA_X1 _2126_ (
  .A(_0924_),
  .B(_0923_),
  .CI(_0890_),
  .CO(_0925_),
  .S(_0926_)
);

FA_X1 _2127_ (
  .A(_0927_),
  .B(_0928_),
  .CI(_0895_),
  .CO(_0929_),
  .S(_0930_)
);

FA_X1 _2128_ (
  .A(_0888_),
  .B(_0930_),
  .CI(_0896_),
  .CO(_0931_),
  .S(_0932_)
);

FA_X1 _2129_ (
  .A(_0926_),
  .B(_0892_),
  .CI(_0932_),
  .CO(_0933_),
  .S(_0934_)
);

FA_X1 _2130_ (
  .A(_0833_),
  .B(_0866_),
  .CI(_0808_),
  .CO(_0935_),
  .S(_0936_)
);

FA_X1 _2131_ (
  .A(_0937_),
  .B(_0938_),
  .CI(_0902_),
  .CO(_0939_),
  .S(_0940_)
);

FA_X1 _2132_ (
  .A(_0898_),
  .B(_0940_),
  .CI(_0906_),
  .CO(_0943_),
  .S(_0944_)
);

FA_X1 _2133_ (
  .A(_0934_),
  .B(_0900_),
  .CI(_0944_),
  .CO(_0945_),
  .S(_0946_)
);

FA_X1 _2134_ (
  .A(_0947_),
  .B(_0948_),
  .CI(_0911_),
  .CO(_0949_),
  .S(_0950_)
);

FA_X1 _2135_ (
  .A(_0951_),
  .B(_0952_),
  .CI(_0953_),
  .CO(_0954_),
  .S(_0955_)
);

FA_X1 _2136_ (
  .A(_0924_),
  .B(_0956_),
  .CI(_0890_),
  .CO(_0957_),
  .S(_0958_)
);

FA_X1 _2137_ (
  .A(_0928_),
  .B(_0959_),
  .CI(_0960_),
  .CO(_0961_),
  .S(_0962_)
);

FA_X1 _2138_ (
  .A(_0922_),
  .B(_0962_),
  .CI(_0929_),
  .CO(_0963_),
  .S(_0964_)
);

FA_X1 _2139_ (
  .A(_0958_),
  .B(_0925_),
  .CI(_0964_),
  .CO(_0965_),
  .S(_0966_)
);

FA_X1 _2140_ (
  .A(_0833_),
  .B(_0866_),
  .CI(_0895_),
  .CO(_0967_),
  .S(_0968_)
);

FA_X1 _2141_ (
  .A(_0969_),
  .B(_0970_),
  .CI(_0935_),
  .CO(_0971_),
  .S(_0972_)
);

FA_X1 _2142_ (
  .A(_0974_),
  .B(_0975_),
  .CI(_0976_),
  .CO(_0977_),
  .S(_0978_)
);

FA_X1 _2143_ (
  .A(_0966_),
  .B(_0933_),
  .CI(_0978_),
  .CO(_0979_),
  .S(_0980_)
);

FA_X1 _2144_ (
  .A(_0981_),
  .B(_0982_),
  .CI(_0983_),
  .CO(_0984_),
  .S(_0985_)
);

FA_X1 _2145_ (
  .A(_0951_),
  .B(_0986_),
  .CI(_0952_),
  .CO(_0987_),
  .S(_0988_)
);

FA_X1 _2146_ (
  .A(_0924_),
  .B(_0989_),
  .CI(_0890_),
  .CO(_0990_),
  .S(_0991_)
);

FA_X1 _2147_ (
  .A(_0992_),
  .B(_0993_),
  .CI(_0960_),
  .CO(_0994_),
  .S(_0995_)
);

FA_X1 _2148_ (
  .A(_0995_),
  .B(_0961_),
  .CI(_0996_),
  .CO(_0997_),
  .S(_0998_)
);

FA_X1 _2149_ (
  .A(_0998_),
  .B(_0991_),
  .CI(_0957_),
  .CO(_0999_),
  .S(_1000_)
);

FA_X1 _2150_ (
  .A(_1001_),
  .B(_1002_),
  .CI(_1003_),
  .CO(_1004_),
  .S(_1005_)
);

FA_X1 _2151_ (
  .A(_1005_),
  .B(_1006_),
  .CI(_0903_),
  .CO(_1007_),
  .S(_1008_)
);

FA_X1 _2152_ (
  .A(_1009_),
  .B(_1008_),
  .CI(_1010_),
  .CO(_1011_),
  .S(_1012_)
);

FA_X1 _2153_ (
  .A(_1000_),
  .B(_0965_),
  .CI(_1012_),
  .CO(_1013_),
  .S(_1014_)
);

FA_X1 _2154_ (
  .A(_1014_),
  .B(_0979_),
  .CI(_1015_),
  .CO(_1016_),
  .S(_1017_)
);

FA_X1 _2155_ (
  .A(_1018_),
  .B(_0984_),
  .CI(_1019_),
  .CO(_1020_),
  .S(_1021_)
);

FA_X1 _2156_ (
  .A(_1022_),
  .B(_1023_),
  .CI(_1024_),
  .CO(_1025_),
  .S(_1026_)
);

FA_X1 _2157_ (
  .A(_1027_),
  .B(_1028_),
  .CI(_0994_),
  .CO(_1029_),
  .S(_1030_)
);

FA_X1 _2158_ (
  .A(_0990_),
  .B(_1030_),
  .CI(_0991_),
  .CO(_1031_),
  .S(_1032_)
);

FA_X1 _2159_ (
  .A(_1001_),
  .B(_1033_),
  .CI(_1003_),
  .CO(_1034_),
  .S(_1035_)
);

FA_X1 _2160_ (
  .A(_1035_),
  .B(_1004_),
  .CI(_0936_),
  .CO(_1036_),
  .S(_1037_)
);

FA_X1 _2161_ (
  .A(_0997_),
  .B(_1038_),
  .CI(_1039_),
  .CO(_1040_),
  .S(_1041_)
);

FA_X1 _2162_ (
  .A(_1032_),
  .B(_0999_),
  .CI(_1041_),
  .CO(_1042_),
  .S(_1043_)
);

FA_X1 _2163_ (
  .A(_1043_),
  .B(_1013_),
  .CI(_1044_),
  .CO(_1045_),
  .S(_1046_)
);

FA_X1 _2164_ (
  .A(_1047_),
  .B(_1048_),
  .CI(_1049_),
  .CO(_1050_),
  .S(_1051_)
);

FA_X1 _2165_ (
  .A(_1052_),
  .B(_1053_),
  .CI(_1054_),
  .CO(_1055_),
  .S(_1056_)
);

FA_X1 _2166_ (
  .A(_1027_),
  .B(_1057_),
  .CI(_1058_),
  .CO(_1059_),
  .S(_1060_)
);

FA_X1 _2167_ (
  .A(_0990_),
  .B(_1060_),
  .CI(_0991_),
  .CO(_1061_),
  .S(_1062_)
);

FA_X1 _2168_ (
  .A(_0993_),
  .B(_0928_),
  .CI(_0960_),
  .CO(_1063_),
  .S(_1064_)
);

FA_X1 _2169_ (
  .A(_1034_),
  .B(_1064_),
  .CI(_0968_),
  .CO(_1065_),
  .S(_1066_)
);

FA_X1 _2170_ (
  .A(_1066_),
  .B(_1036_),
  .CI(_1067_),
  .CO(_1068_),
  .S(_1069_)
);

FA_X1 _2171_ (
  .A(_1069_),
  .B(_1062_),
  .CI(_1031_),
  .CO(_1070_),
  .S(_1071_)
);

FA_X1 _2172_ (
  .A(_0973_),
  .B(_0875_),
  .CI(_1072_),
  .CO(_1073_),
  .S(_1074_)
);

FA_X1 _2173_ (
  .A(_1075_),
  .B(_1076_),
  .CI(_1077_),
  .CO(_1078_),
  .S(_1079_)
);

FA_X1 _2174_ (
  .A(_1071_),
  .B(_1042_),
  .CI(_1080_),
  .CO(_1081_),
  .S(_1082_)
);

FA_X1 _2175_ (
  .A(_1083_),
  .B(_1084_),
  .CI(_1085_),
  .CO(_1086_),
  .S(_1087_)
);

HA_X1 _2176_ (
  .A(result[0]),
  .B(\ext_mult_res[0] ),
  .CO(_1088_),
  .S(_1089_)
);

HA_X1 _2177_ (
  .A(result[1]),
  .B(\ext_mult_res[1] ),
  .CO(_1090_),
  .S(_1091_)
);

HA_X1 _2178_ (
  .A(result[2]),
  .B(\ext_mult_res[2] ),
  .CO(_1092_),
  .S(_1093_)
);

HA_X1 _2179_ (
  .A(result[3]),
  .B(\ext_mult_res[3] ),
  .CO(_1094_),
  .S(_1095_)
);

HA_X1 _2180_ (
  .A(result[4]),
  .B(\ext_mult_res[4] ),
  .CO(_1096_),
  .S(_1097_)
);

HA_X1 _2181_ (
  .A(result[5]),
  .B(\ext_mult_res[5] ),
  .CO(_1098_),
  .S(_1099_)
);

HA_X1 _2182_ (
  .A(result[6]),
  .B(\ext_mult_res[6] ),
  .CO(_1100_),
  .S(_1101_)
);

HA_X1 _2183_ (
  .A(result[7]),
  .B(\ext_mult_res[7] ),
  .CO(_1102_),
  .S(_1103_)
);

HA_X1 _2184_ (
  .A(result[8]),
  .B(\ext_mult_res[8] ),
  .CO(_1104_),
  .S(_1105_)
);

HA_X1 _2185_ (
  .A(result[9]),
  .B(\ext_mult_res[9] ),
  .CO(_1106_),
  .S(_1107_)
);

HA_X1 _2186_ (
  .A(result[10]),
  .B(\ext_mult_res[10] ),
  .CO(_1108_),
  .S(_1109_)
);

HA_X1 _2187_ (
  .A(result[11]),
  .B(\ext_mult_res[11] ),
  .CO(_1110_),
  .S(_1111_)
);

HA_X1 _2188_ (
  .A(result[12]),
  .B(\ext_mult_res[12] ),
  .CO(_1112_),
  .S(_1113_)
);

HA_X1 _2189_ (
  .A(result[13]),
  .B(\ext_mult_res[13] ),
  .CO(_1114_),
  .S(_1115_)
);

HA_X1 _2190_ (
  .A(result[14]),
  .B(\ext_mult_res[14] ),
  .CO(_1116_),
  .S(_1117_)
);

HA_X1 _2191_ (
  .A(result[15]),
  .B(\ext_mult_res[15] ),
  .CO(_1118_),
  .S(_1119_)
);

HA_X1 _2192_ (
  .A(result[16]),
  .B(\ext_mult_res[16] ),
  .CO(_1120_),
  .S(_1121_)
);

HA_X1 _2193_ (
  .A(result[17]),
  .B(\ext_mult_res[17] ),
  .CO(_1122_),
  .S(_1123_)
);

HA_X1 _2194_ (
  .A(result[18]),
  .B(\ext_mult_res[18] ),
  .CO(_1124_),
  .S(_1125_)
);

HA_X1 _2195_ (
  .A(result[19]),
  .B(\ext_mult_res[18] ),
  .CO(_1126_),
  .S(_1127_)
);

HA_X1 _2196_ (
  .A(result[20]),
  .B(\ext_mult_res[18] ),
  .CO(_1128_),
  .S(_1129_)
);

HA_X1 _2197_ (
  .A(_1130_),
  .B(_1131_),
  .CO(_1132_),
  .S(_1133_)
);

HA_X1 _2198_ (
  .A(_0685_),
  .B(_1132_),
  .CO(_1134_),
  .S(_1135_)
);

HA_X1 _2199_ (
  .A(_0693_),
  .B(_1134_),
  .CO(_1136_),
  .S(_1137_)
);

HA_X1 _2200_ (
  .A(_1138_),
  .B(_1139_),
  .CO(_0717_),
  .S(_1140_)
);

HA_X1 _2201_ (
  .A(_1141_),
  .B(_0692_),
  .CO(_1142_),
  .S(_1143_)
);

HA_X1 _2202_ (
  .A(_1143_),
  .B(_1136_),
  .CO(_1144_),
  .S(_1145_)
);

HA_X1 _2203_ (
  .A(_0719_),
  .B(_1142_),
  .CO(_1146_),
  .S(_1147_)
);

HA_X1 _2204_ (
  .A(_1147_),
  .B(_1144_),
  .CO(_1148_),
  .S(_1149_)
);

HA_X1 _2205_ (
  .A(_1150_),
  .B(_1151_),
  .CO(_1152_),
  .S(_1153_)
);

HA_X1 _2206_ (
  .A(_1154_),
  .B(_0718_),
  .CO(_1155_),
  .S(_1156_)
);

HA_X1 _2207_ (
  .A(_1156_),
  .B(_1146_),
  .CO(_1157_),
  .S(_1158_)
);

HA_X1 _2208_ (
  .A(_1158_),
  .B(_1148_),
  .CO(_1159_),
  .S(_1160_)
);

HA_X1 _2209_ (
  .A(_0764_),
  .B(_1161_),
  .CO(_0767_),
  .S(_1162_)
);

HA_X1 _2210_ (
  .A(_1163_),
  .B(_1162_),
  .CO(_0780_),
  .S(_1164_)
);

HA_X1 _2211_ (
  .A(_0782_),
  .B(_1165_),
  .CO(_1166_),
  .S(_1167_)
);

HA_X1 _2212_ (
  .A(_1167_),
  .B(_1168_),
  .CO(_1169_),
  .S(_1170_)
);

HA_X1 _2213_ (
  .A(_1171_),
  .B(_1155_),
  .CO(_1168_),
  .S(_1172_)
);

HA_X1 _2214_ (
  .A(_1170_),
  .B(_1173_),
  .CO(_1174_),
  .S(_1175_)
);

HA_X1 _2215_ (
  .A(_1172_),
  .B(_1157_),
  .CO(_1173_),
  .S(_1176_)
);

HA_X1 _2216_ (
  .A(_0764_),
  .B(_0768_),
  .CO(_0847_),
  .S(_1178_)
);

HA_X1 _2217_ (
  .A(_1179_),
  .B(_0781_),
  .CO(_1180_),
  .S(_1181_)
);

HA_X1 _2218_ (
  .A(_1181_),
  .B(_1166_),
  .CO(_1182_),
  .S(_1183_)
);

HA_X1 _2219_ (
  .A(_1183_),
  .B(_1169_),
  .CO(_1184_),
  .S(_1185_)
);

HA_X1 _2220_ (
  .A(_0763_),
  .B(_0764_),
  .CO(_1072_),
  .S(_0941_)
);

HA_X1 _2221_ (
  .A(_0814_),
  .B(_0941_),
  .CO(_1186_),
  .S(_1187_)
);

HA_X1 _2222_ (
  .A(_0851_),
  .B(_1180_),
  .CO(_1188_),
  .S(_1189_)
);

HA_X1 _2223_ (
  .A(_1189_),
  .B(_1182_),
  .CO(_1190_),
  .S(_1191_)
);

HA_X1 _2224_ (
  .A(_0875_),
  .B(_1072_),
  .CO(_0910_),
  .S(_1192_)
);

HA_X1 _2225_ (
  .A(_0840_),
  .B(_1192_),
  .CO(_1193_),
  .S(_1194_)
);

HA_X1 _2226_ (
  .A(_0881_),
  .B(_0850_),
  .CO(_1195_),
  .S(_1196_)
);

HA_X1 _2227_ (
  .A(_1196_),
  .B(_1188_),
  .CO(_1197_),
  .S(_1198_)
);

HA_X1 _2228_ (
  .A(_1199_),
  .B(_0918_),
  .CO(_1200_),
  .S(_1201_)
);

HA_X1 _2229_ (
  .A(_1195_),
  .B(_1201_),
  .CO(_1202_),
  .S(_1203_)
);

HA_X1 _2230_ (
  .A(_1204_),
  .B(_1205_),
  .CO(_1206_),
  .S(_1207_)
);

HA_X1 _2231_ (
  .A(_1207_),
  .B(_1200_),
  .CO(_1208_),
  .S(_1209_)
);

HA_X1 _2232_ (
  .A(_1210_),
  .B(_1072_),
  .CO(_1019_),
  .S(_0981_)
);

HA_X1 _2233_ (
  .A(_1211_),
  .B(_0949_),
  .CO(_1212_),
  .S(_1213_)
);

HA_X1 _2234_ (
  .A(_1213_),
  .B(_1206_),
  .CO(_1214_),
  .S(_1215_)
);

HA_X1 _2235_ (
  .A(_0764_),
  .B(_0874_),
  .CO(_1217_),
  .S(_1218_)
);

HA_X1 _2236_ (
  .A(_0977_),
  .B(_1218_),
  .CO(_1049_),
  .S(_1219_)
);

HA_X1 _2237_ (
  .A(_1021_),
  .B(_1212_),
  .CO(_1220_),
  .S(_1221_)
);

HA_X1 _2238_ (
  .A(_1222_),
  .B(_1216_),
  .CO(_1223_),
  .S(_1224_)
);

HA_X1 _2239_ (
  .A(_0941_),
  .B(_0942_),
  .CO(_1225_),
  .S(_1226_)
);

HA_X1 _2240_ (
  .A(_1226_),
  .B(_1217_),
  .CO(_1077_),
  .S(_1227_)
);

HA_X1 _2241_ (
  .A(_1011_),
  .B(_1227_),
  .CO(_1085_),
  .S(_1228_)
);

HA_X1 _2242_ (
  .A(_1051_),
  .B(_1020_),
  .CO(_1229_),
  .S(_1230_)
);

HA_X1 _2243_ (
  .A(_1074_),
  .B(_1225_),
  .CO(_1231_),
  .S(_1076_)
);

HA_X1 _2244_ (
  .A(_1087_),
  .B(_1050_),
  .CO(_1232_),
  .S(_1233_)
);

HA_X1 _2245_ (
  .A(_1176_),
  .B(_1159_),
  .CO(_1177_),
  .S(_1234_)
);

DFF_X1 \ext_mult_res[0]$_DFFE_PP_  (
  .D(_0000_),
  .CK(clk),
  .Q(\ext_mult_res[0] ),
  .QN(_0675_)
);

DFF_X1 \ext_mult_res[10]$_DFFE_PP_  (
  .D(_0010_),
  .CK(clk),
  .Q(\ext_mult_res[10] ),
  .QN(_0666_)
);

DFF_X1 \ext_mult_res[11]$_DFFE_PP_  (
  .D(_0011_),
  .CK(clk),
  .Q(\ext_mult_res[11] ),
  .QN(_0665_)
);

DFF_X1 \ext_mult_res[12]$_DFFE_PP_  (
  .D(_0012_),
  .CK(clk),
  .Q(\ext_mult_res[12] ),
  .QN(_0664_)
);

DFF_X1 \ext_mult_res[13]$_DFFE_PP_  (
  .D(_0013_),
  .CK(clk),
  .Q(\ext_mult_res[13] ),
  .QN(_0663_)
);

DFF_X1 \ext_mult_res[14]$_DFFE_PP_  (
  .D(_0014_),
  .CK(clk),
  .Q(\ext_mult_res[14] ),
  .QN(_0662_)
);

DFF_X1 \ext_mult_res[15]$_DFFE_PP_  (
  .D(_0015_),
  .CK(clk),
  .Q(\ext_mult_res[15] ),
  .QN(_0661_)
);

DFF_X1 \ext_mult_res[16]$_DFFE_PP_  (
  .D(_0016_),
  .CK(clk),
  .Q(\ext_mult_res[16] ),
  .QN(_0660_)
);

DFF_X1 \ext_mult_res[17]$_DFFE_PP_  (
  .D(_0017_),
  .CK(clk),
  .Q(\ext_mult_res[17] ),
  .QN(_0659_)
);

DFF_X1 \ext_mult_res[1]$_DFFE_PP_  (
  .D(_0001_),
  .CK(clk),
  .Q(\ext_mult_res[1] ),
  .QN(_0677_)
);

DFF_X1 \ext_mult_res[21]$_DFFE_PP_  (
  .D(_0018_),
  .CK(clk),
  .Q(\ext_mult_res[18] ),
  .QN(_0658_)
);

DFF_X1 \ext_mult_res[2]$_DFFE_PP_  (
  .D(_0002_),
  .CK(clk),
  .Q(\ext_mult_res[2] ),
  .QN(_0674_)
);

DFF_X1 \ext_mult_res[3]$_DFFE_PP_  (
  .D(_0003_),
  .CK(clk),
  .Q(\ext_mult_res[3] ),
  .QN(_0673_)
);

DFF_X1 \ext_mult_res[4]$_DFFE_PP_  (
  .D(_0004_),
  .CK(clk),
  .Q(\ext_mult_res[4] ),
  .QN(_0672_)
);

DFF_X1 \ext_mult_res[5]$_DFFE_PP_  (
  .D(_0005_),
  .CK(clk),
  .Q(\ext_mult_res[5] ),
  .QN(_0671_)
);

DFF_X1 \ext_mult_res[6]$_DFFE_PP_  (
  .D(_0006_),
  .CK(clk),
  .Q(\ext_mult_res[6] ),
  .QN(_0670_)
);

DFF_X1 \ext_mult_res[7]$_DFFE_PP_  (
  .D(_0007_),
  .CK(clk),
  .Q(\ext_mult_res[7] ),
  .QN(_0669_)
);

DFF_X1 \ext_mult_res[8]$_DFFE_PP_  (
  .D(_0008_),
  .CK(clk),
  .Q(\ext_mult_res[8] ),
  .QN(_0668_)
);

DFF_X1 \ext_mult_res[9]$_DFFE_PP_  (
  .D(_0009_),
  .CK(clk),
  .Q(\ext_mult_res[9] ),
  .QN(_0667_)
);

DFF_X1 \result[0]$_DFFE_PP_  (
  .D(_0019_),
  .CK(clk),
  .Q(result[0]),
  .QN(_0657_)
);

DFF_X1 \result[10]$_DFFE_PP_  (
  .D(_0029_),
  .CK(clk),
  .Q(result[10]),
  .QN(_0648_)
);

DFF_X1 \result[11]$_DFFE_PP_  (
  .D(_0030_),
  .CK(clk),
  .Q(result[11]),
  .QN(_0647_)
);

DFF_X1 \result[12]$_DFFE_PP_  (
  .D(_0031_),
  .CK(clk),
  .Q(result[12]),
  .QN(_0646_)
);

DFF_X1 \result[13]$_DFFE_PP_  (
  .D(_0032_),
  .CK(clk),
  .Q(result[13]),
  .QN(_0645_)
);

DFF_X1 \result[14]$_DFFE_PP_  (
  .D(_0033_),
  .CK(clk),
  .Q(result[14]),
  .QN(_0644_)
);

DFF_X1 \result[15]$_DFFE_PP_  (
  .D(_0034_),
  .CK(clk),
  .Q(result[15]),
  .QN(_0643_)
);

DFF_X1 \result[16]$_DFFE_PP_  (
  .D(_0035_),
  .CK(clk),
  .Q(result[16]),
  .QN(_0642_)
);

DFF_X1 \result[17]$_DFFE_PP_  (
  .D(_0036_),
  .CK(clk),
  .Q(result[17]),
  .QN(_0641_)
);

DFF_X1 \result[18]$_DFFE_PP_  (
  .D(_0037_),
  .CK(clk),
  .Q(result[18]),
  .QN(_0640_)
);

DFF_X1 \result[19]$_DFFE_PP_  (
  .D(_0038_),
  .CK(clk),
  .Q(result[19]),
  .QN(_0639_)
);

DFF_X1 \result[1]$_DFFE_PP_  (
  .D(_0020_),
  .CK(clk),
  .Q(result[1]),
  .QN(_0676_)
);

DFF_X1 \result[20]$_DFFE_PP_  (
  .D(_0039_),
  .CK(clk),
  .Q(result[20]),
  .QN(_0638_)
);

DFF_X1 \result[21]$_DFFE_PP_  (
  .D(_0040_),
  .CK(clk),
  .Q(result[21]),
  .QN(_0637_)
);

DFF_X1 \result[2]$_DFFE_PP_  (
  .D(_0021_),
  .CK(clk),
  .Q(result[2]),
  .QN(_0656_)
);

DFF_X1 \result[3]$_DFFE_PP_  (
  .D(_0022_),
  .CK(clk),
  .Q(result[3]),
  .QN(_0655_)
);

DFF_X1 \result[4]$_DFFE_PP_  (
  .D(_0023_),
  .CK(clk),
  .Q(result[4]),
  .QN(_0654_)
);

DFF_X1 \result[5]$_DFFE_PP_  (
  .D(_0024_),
  .CK(clk),
  .Q(result[5]),
  .QN(_0653_)
);

DFF_X1 \result[6]$_DFFE_PP_  (
  .D(_0025_),
  .CK(clk),
  .Q(result[6]),
  .QN(_0652_)
);

DFF_X1 \result[7]$_DFFE_PP_  (
  .D(_0026_),
  .CK(clk),
  .Q(result[7]),
  .QN(_0651_)
);

DFF_X1 \result[8]$_DFFE_PP_  (
  .D(_0027_),
  .CK(clk),
  .Q(result[8]),
  .QN(_0650_)
);

DFF_X1 \result[9]$_DFFE_PP_  (
  .D(_0028_),
  .CK(clk),
  .Q(result[9]),
  .QN(_0649_)
);
endmodule //$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac

module \$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 (input clk,
 input ena, input dclr, input [7:0] din, input [10:0] coef, output [21:0] result);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire _0032_;
wire _0033_;
wire _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire _0066_;
wire _0067_;
wire _0068_;
wire _0069_;
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0333_;
wire _0339_;
wire _0341_;
wire _0348_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0367_;
wire _0368_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
wire _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
wire _0444_;
wire _0445_;
wire _0446_;
wire _0447_;
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire _0658_;
wire _0659_;
wire _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire _0673_;
wire _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire _0679_;
wire _0680_;
wire _0684_;
wire _0685_;
wire _0689_;
wire _0690_;
wire _0692_;
wire _0693_;
wire _0697_;
wire _0698_;
wire _0699_;
wire _0700_;
wire _0701_;
wire _0702_;
wire _0706_;
wire _0707_;
wire _0711_;
wire _0712_;
wire _0713_;
wire _0714_;
wire _0715_;
wire _0716_;
wire _0717_;
wire _0718_;
wire _0719_;
wire _0723_;
wire _0724_;
wire _0728_;
wire _0729_;
wire _0730_;
wire _0731_;
wire _0732_;
wire _0733_;
wire _0734_;
wire _0735_;
wire _0738_;
wire _0739_;
wire _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0751_;
wire _0752_;
wire _0756_;
wire _0757_;
wire _0761_;
wire _0762_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire _0780_;
wire _0781_;
wire _0782_;
wire _0783_;
wire _0784_;
wire _0785_;
wire _0786_;
wire _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire _0795_;
wire _0796_;
wire _0798_;
wire _0799_;
wire _0803_;
wire _0804_;
wire _0805_;
wire _0806_;
wire _0809_;
wire _0810_;
wire _0811_;
wire _0812_;
wire _0813_;
wire _0814_;
wire _0815_;
wire _0816_;
wire _0817_;
wire _0818_;
wire _0819_;
wire _0820_;
wire _0821_;
wire _0822_;
wire _0823_;
wire _0824_;
wire _0825_;
wire _0829_;
wire _0830_;
wire _0831_;
wire _0832_;
wire _0835_;
wire _0836_;
wire _0837_;
wire _0838_;
wire _0839_;
wire _0840_;
wire _0841_;
wire _0842_;
wire _0843_;
wire _0844_;
wire _0845_;
wire _0846_;
wire _0847_;
wire _0848_;
wire _0849_;
wire _0850_;
wire _0851_;
wire _0852_;
wire _0853_;
wire _0854_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0860_;
wire _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0867_;
wire _0868_;
wire _0869_;
wire _0870_;
wire _0871_;
wire _0872_;
wire _0874_;
wire _0875_;
wire _0876_;
wire _0877_;
wire _0878_;
wire _0879_;
wire _0880_;
wire _0881_;
wire _0882_;
wire _0883_;
wire _0884_;
wire _0885_;
wire _0886_;
wire _0888_;
wire _0889_;
wire _0890_;
wire _0891_;
wire _0892_;
wire _0893_;
wire _0896_;
wire _0897_;
wire _0898_;
wire _0899_;
wire _0900_;
wire _0901_;
wire _0902_;
wire _0903_;
wire _0904_;
wire _0905_;
wire _0906_;
wire _0907_;
wire _0908_;
wire _0909_;
wire _0910_;
wire _0911_;
wire _0912_;
wire _0913_;
wire _0914_;
wire _0915_;
wire _0916_;
wire _0917_;
wire _0918_;
wire _0919_;
wire _0920_;
wire _0921_;
wire _0922_;
wire _0923_;
wire _0924_;
wire _0925_;
wire _0926_;
wire _0929_;
wire _0930_;
wire _0931_;
wire _0932_;
wire _0933_;
wire _0934_;
wire _0935_;
wire _0936_;
wire _0937_;
wire _0938_;
wire _0939_;
wire _0940_;
wire _0941_;
wire _0942_;
wire _0943_;
wire _0944_;
wire _0945_;
wire _0946_;
wire _0947_;
wire _0948_;
wire _0949_;
wire _0950_;
wire _0951_;
wire _0952_;
wire _0953_;
wire _0954_;
wire _0955_;
wire _0956_;
wire _0957_;
wire _0958_;
wire _0959_;
wire _0961_;
wire _0962_;
wire _0963_;
wire _0964_;
wire _0965_;
wire _0966_;
wire _0967_;
wire _0968_;
wire _0969_;
wire _0970_;
wire _0971_;
wire _0972_;
wire _0973_;
wire _0974_;
wire _0975_;
wire _0976_;
wire _0977_;
wire _0978_;
wire _0979_;
wire _0980_;
wire _0981_;
wire _0982_;
wire _0983_;
wire _0984_;
wire _0985_;
wire _0986_;
wire _0987_;
wire _0988_;
wire _0989_;
wire _0990_;
wire _0991_;
wire _0992_;
wire _0993_;
wire _0994_;
wire _0995_;
wire _0996_;
wire _0997_;
wire _0998_;
wire _0999_;
wire _1000_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire \ext_mult_res[0] ;
wire \ext_mult_res[10] ;
wire \ext_mult_res[11] ;
wire \ext_mult_res[12] ;
wire \ext_mult_res[13] ;
wire \ext_mult_res[14] ;
wire \ext_mult_res[15] ;
wire \ext_mult_res[16] ;
wire \ext_mult_res[17] ;
wire \ext_mult_res[18] ;
wire \ext_mult_res[1] ;
wire \ext_mult_res[2] ;
wire \ext_mult_res[3] ;
wire \ext_mult_res[4] ;
wire \ext_mult_res[5] ;
wire \ext_mult_res[6] ;
wire \ext_mult_res[7] ;
wire \ext_mult_res[8] ;
wire \ext_mult_res[9] ;
wire \logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ;
wire \logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ;

BUF_X1 _1235_ (
  .A(din[0]),
  .Z(_0326_)
);

BUF_X1 _1245_ (
  .A(din[1]),
  .Z(_0333_)
);

BUF_X1 _1255_ (
  .A(din[2]),
  .Z(_0339_)
);

BUF_X1 _1258_ (
  .A(din[3]),
  .Z(_0341_)
);

BUF_X1 _1279_ (
  .A(din[6]),
  .Z(_0348_)
);

BUF_X1 _1292_ (
  .A(din[4]),
  .Z(_0354_)
);

BUF_X1 _1294_ (
  .A(din[5]),
  .Z(_0355_)
);

BUF_X8 _1299_ (
  .A(din[7]),
  .Z(_0356_)
);

BUF_X4 _1306_ (
  .A(coef[9]),
  .Z(_0358_)
);

NAND2_X1 _1307_ (
  .A1(_0326_),
  .A2(_0358_),
  .ZN(_0795_)
);

BUF_X4 _1316_ (
  .A(coef[10]),
  .Z(_0359_)
);

NAND2_X1 _1317_ (
  .A1(_0326_),
  .A2(_0359_),
  .ZN(_0821_)
);

INV_X1 _1318_ (
  .A(_0821_),
  .ZN(_0854_)
);

NAND2_X1 _1324_ (
  .A1(_0333_),
  .A2(_0359_),
  .ZN(_0360_)
);

INV_X1 _1325_ (
  .A(_0360_),
  .ZN(_0852_)
);

NAND2_X1 _1326_ (
  .A1(_0339_),
  .A2(_0358_),
  .ZN(_0361_)
);

INV_X1 _1327_ (
  .A(_0361_),
  .ZN(_0853_)
);

NAND2_X1 _1334_ (
  .A1(_0339_),
  .A2(_0359_),
  .ZN(_0362_)
);

INV_X1 _1335_ (
  .A(_0362_),
  .ZN(_0882_)
);

NAND2_X1 _1336_ (
  .A1(_0341_),
  .A2(_0358_),
  .ZN(_0885_)
);

INV_X1 _1342_ (
  .A(_1177_),
  .ZN(_0792_)
);

NAND2_X1 _1343_ (
  .A1(din[3]),
  .A2(_0359_),
  .ZN(_0919_)
);

INV_X1 _1344_ (
  .A(_0919_),
  .ZN(_0951_)
);

NAND2_X1 _1349_ (
  .A1(_0354_),
  .A2(_0359_),
  .ZN(_0363_)
);

INV_X1 _1350_ (
  .A(_0363_),
  .ZN(_0952_)
);

NAND2_X1 _1351_ (
  .A1(din[5]),
  .A2(_0358_),
  .ZN(_0364_)
);

INV_X1 _1352_ (
  .A(_0364_),
  .ZN(_0953_)
);

NAND2_X1 _1356_ (
  .A1(_0355_),
  .A2(_0359_),
  .ZN(_0365_)
);

INV_X1 _1357_ (
  .A(_0365_),
  .ZN(_0986_)
);

NAND2_X1 _1358_ (
  .A1(_0348_),
  .A2(_0358_),
  .ZN(_0992_)
);

INV_X1 _1360_ (
  .A(_0993_),
  .ZN(_1022_)
);

NAND2_X2 _1361_ (
  .A1(din[6]),
  .A2(_0359_),
  .ZN(_1052_)
);

INV_X2 _1362_ (
  .A(_1052_),
  .ZN(_1023_)
);

NAND2_X2 _1363_ (
  .A1(_0356_),
  .A2(_0358_),
  .ZN(_1053_)
);

INV_X4 _1364_ (
  .A(_1053_),
  .ZN(_1024_)
);

INV_X1 _1365_ (
  .A(_0987_),
  .ZN(_1027_)
);

INV_X1 _1366_ (
  .A(_0874_),
  .ZN(_0905_)
);

INV_X1 _1368_ (
  .A(_0785_),
  .ZN(_0786_)
);

INV_X1 _1370_ (
  .A(_0875_),
  .ZN(_0969_)
);

NAND2_X1 _1373_ (
  .A1(_0333_),
  .A2(_0358_),
  .ZN(_0822_)
);

INV_X1 _1374_ (
  .A(_0903_),
  .ZN(_0904_)
);

NAND2_X1 _1375_ (
  .A1(_0354_),
  .A2(_0358_),
  .ZN(_0920_)
);

INV_X1 _1376_ (
  .A(_0936_),
  .ZN(_0938_)
);

INV_X1 _1377_ (
  .A(_0968_),
  .ZN(_0970_)
);

INV_X1 _1378_ (
  .A(_1088_),
  .ZN(_0678_)
);

INV_X1 _1381_ (
  .A(_1152_),
  .ZN(_0787_)
);

INV_X1 _1382_ (
  .A(_1186_),
  .ZN(_0879_)
);

INV_X1 _1383_ (
  .A(_1193_),
  .ZN(_0916_)
);

NAND2_X1 _1384_ (
  .A1(_0356_),
  .A2(_0359_),
  .ZN(_1054_)
);

INV_X1 _1385_ (
  .A(_1029_),
  .ZN(_1067_)
);

INV_X1 _1386_ (
  .A(_0752_),
  .ZN(_0775_)
);

INV_X1 _1387_ (
  .A(_0769_),
  .ZN(_0771_)
);

INV_X1 _1388_ (
  .A(_0856_),
  .ZN(_0862_)
);

INV_X1 _1389_ (
  .A(_0884_),
  .ZN(_0890_)
);

INV_X1 _1390_ (
  .A(_0912_),
  .ZN(_0913_)
);

INV_X1 _1391_ (
  .A(_0950_),
  .ZN(_1204_)
);

INV_X1 _1392_ (
  .A(_0955_),
  .ZN(_0956_)
);

INV_X1 _1393_ (
  .A(_0985_),
  .ZN(_1211_)
);

INV_X1 _1394_ (
  .A(_0988_),
  .ZN(_0989_)
);

INV_X1 _1395_ (
  .A(_1026_),
  .ZN(_1028_)
);

INV_X1 _1396_ (
  .A(_1037_),
  .ZN(_1038_)
);

INV_X1 _1397_ (
  .A(_1056_),
  .ZN(_1057_)
);

INV_X1 _1398_ (
  .A(_1079_),
  .ZN(_1080_)
);

INV_X1 _1399_ (
  .A(_0689_),
  .ZN(_0699_)
);

INV_X1 _1400_ (
  .A(_0751_),
  .ZN(_0745_)
);

INV_X1 _1401_ (
  .A(_0776_),
  .ZN(_0770_)
);

INV_X1 _1402_ (
  .A(_0855_),
  .ZN(_0891_)
);

INV_X1 _1403_ (
  .A(_0883_),
  .ZN(_0924_)
);

INV_X1 _1404_ (
  .A(_0954_),
  .ZN(_0996_)
);

INV_X1 _1405_ (
  .A(_1007_),
  .ZN(_1039_)
);

INV_X1 _1406_ (
  .A(_1025_),
  .ZN(_1058_)
);

INV_X1 _1407_ (
  .A(_0702_),
  .ZN(_1141_)
);

INV_X1 _1408_ (
  .A(_0714_),
  .ZN(_0715_)
);

INV_X1 _1409_ (
  .A(_0711_),
  .ZN(_1150_)
);

INV_X1 _1410_ (
  .A(_0734_),
  .ZN(_1154_)
);

INV_X1 _1413_ (
  .A(_0723_),
  .ZN(_0774_)
);

INV_X1 _1414_ (
  .A(_0756_),
  .ZN(_0765_)
);

INV_X1 _1415_ (
  .A(_0728_),
  .ZN(_1163_)
);

INV_X1 _1416_ (
  .A(_0773_),
  .ZN(_0778_)
);

INV_X1 _1417_ (
  .A(_0789_),
  .ZN(_1171_)
);

INV_X1 _1418_ (
  .A(_0743_),
  .ZN(_0811_)
);

INV_X1 _1419_ (
  .A(_0820_),
  .ZN(_1179_)
);

INV_X1 _1420_ (
  .A(_0836_),
  .ZN(_0838_)
);

INV_X1 _1421_ (
  .A(_0809_),
  .ZN(_0837_)
);

INV_X1 _1422_ (
  .A(_0846_),
  .ZN(_0848_)
);

INV_X1 _1423_ (
  .A(_0869_),
  .ZN(_0908_)
);

INV_X1 _1424_ (
  .A(_0880_),
  .ZN(_1199_)
);

INV_X1 _1425_ (
  .A(_0946_),
  .ZN(_0947_)
);

INV_X1 _1426_ (
  .A(_0931_),
  .ZN(_0974_)
);

INV_X1 _1427_ (
  .A(_0945_),
  .ZN(_0982_)
);

INV_X1 _1428_ (
  .A(_0943_),
  .ZN(_1210_)
);

INV_X1 _1429_ (
  .A(_0991_),
  .ZN(_1216_)
);

INV_X1 _1430_ (
  .A(_0963_),
  .ZN(_1009_)
);

INV_X1 _1431_ (
  .A(_1017_),
  .ZN(_1018_)
);

INV_X1 _1432_ (
  .A(_0990_),
  .ZN(_1222_)
);

INV_X1 _1433_ (
  .A(_1046_),
  .ZN(_1047_)
);

INV_X1 _1434_ (
  .A(_1040_),
  .ZN(_1075_)
);

INV_X1 _1435_ (
  .A(_1082_),
  .ZN(_1083_)
);

INV_X1 _1436_ (
  .A(_0701_),
  .ZN(_0716_)
);

INV_X1 _1437_ (
  .A(_0762_),
  .ZN(_0766_)
);

INV_X1 _1438_ (
  .A(_0783_),
  .ZN(_0779_)
);

INV_X1 _1439_ (
  .A(_0788_),
  .ZN(_1165_)
);

INV_X1 _1440_ (
  .A(_0810_),
  .ZN(_0812_)
);

INV_X1 _1441_ (
  .A(_0761_),
  .ZN(_0813_)
);

INV_X1 _1442_ (
  .A(_0803_),
  .ZN(_0839_)
);

INV_X1 _1443_ (
  .A(_0819_),
  .ZN(_0849_)
);

INV_X1 _1444_ (
  .A(_0907_),
  .ZN(_0909_)
);

INV_X1 _1445_ (
  .A(_0914_),
  .ZN(_0948_)
);

INV_X1 _1446_ (
  .A(_0917_),
  .ZN(_1205_)
);

INV_X1 _1447_ (
  .A(_0935_),
  .ZN(_0973_)
);

INV_X1 _1448_ (
  .A(_0972_),
  .ZN(_0975_)
);

INV_X1 _1449_ (
  .A(_0939_),
  .ZN(_0976_)
);

INV_X1 _1450_ (
  .A(_0980_),
  .ZN(_0983_)
);

INV_X1 _1451_ (
  .A(_0967_),
  .ZN(_1006_)
);

INV_X1 _1452_ (
  .A(_0971_),
  .ZN(_1010_)
);

INV_X1 _1453_ (
  .A(_0902_),
  .ZN(_0942_)
);

INV_X1 _1454_ (
  .A(_1016_),
  .ZN(_1048_)
);

INV_X1 _1455_ (
  .A(_1045_),
  .ZN(_1084_)
);

INV_X1 _1456_ (
  .A(_1153_),
  .ZN(_0732_)
);

INV_X1 _1457_ (
  .A(_1170_),
  .ZN(_0790_)
);

INV_X1 _1458_ (
  .A(_1178_),
  .ZN(_0818_)
);

INV_X1 _1459_ (
  .A(_1187_),
  .ZN(_0844_)
);

INV_X1 _1460_ (
  .A(_1194_),
  .ZN(_0876_)
);

INV_X1 _1461_ (
  .A(_1219_),
  .ZN(_1015_)
);

INV_X1 _1462_ (
  .A(_1228_),
  .ZN(_1044_)
);

INV_X1 _1463_ (
  .A(_1140_),
  .ZN(_0700_)
);

INV_X1 _1464_ (
  .A(_1164_),
  .ZN(_0784_)
);

INV_X1 _1465_ (
  .A(_0941_),
  .ZN(_0937_)
);

INV_X1 _1466_ (
  .A(_1173_),
  .ZN(_0791_)
);

BUF_X1 _1467_ (
  .A(ena),
  .Z(_0367_)
);

BUF_X1 _1468_ (
  .A(_0367_),
  .Z(_0368_)
);

INV_X1 _1470_ (
  .A(\ext_mult_res[0] ),
  .ZN(_0370_)
);

BUF_X1 _1471_ (
  .A(_0367_),
  .Z(_0371_)
);

BUF_X1 _1472_ (
  .A(_0371_),
  .Z(_0372_)
);

BUF_X1 _1474_ (
  .A(_0367_),
  .Z(_0373_)
);

MUX2_X1 _1475_ (
  .A(\ext_mult_res[1] ),
  .B(_1133_),
  .S(_0373_),
  .Z(_0001_)
);

BUF_X4 _1476_ (
  .A(_0371_),
  .Z(_0374_)
);

NAND2_X1 _1477_ (
  .A1(_0374_),
  .A2(_1135_),
  .ZN(_0375_)
);

INV_X1 _1478_ (
  .A(\ext_mult_res[2] ),
  .ZN(_0376_)
);

OAI21_X1 _1479_ (
  .A(_0375_),
  .B1(_0376_),
  .B2(_0372_),
  .ZN(_0002_)
);

NAND2_X1 _1480_ (
  .A1(_0374_),
  .A2(_1137_),
  .ZN(_0377_)
);

INV_X1 _1481_ (
  .A(\ext_mult_res[3] ),
  .ZN(_0378_)
);

OAI21_X1 _1482_ (
  .A(_0377_),
  .B1(_0378_),
  .B2(_0372_),
  .ZN(_0003_)
);

NAND2_X1 _1483_ (
  .A1(_0374_),
  .A2(_1145_),
  .ZN(_0379_)
);

INV_X1 _1484_ (
  .A(\ext_mult_res[4] ),
  .ZN(_0380_)
);

OAI21_X1 _1485_ (
  .A(_0379_),
  .B1(_0380_),
  .B2(_0372_),
  .ZN(_0004_)
);

MUX2_X1 _1486_ (
  .A(\ext_mult_res[5] ),
  .B(_1149_),
  .S(_0373_),
  .Z(_0005_)
);

NAND2_X1 _1487_ (
  .A1(_0372_),
  .A2(_1160_),
  .ZN(_0381_)
);

INV_X1 _1488_ (
  .A(\ext_mult_res[6] ),
  .ZN(_0382_)
);

OAI21_X1 _1489_ (
  .A(_0381_),
  .B1(_0382_),
  .B2(_0372_),
  .ZN(_0006_)
);

NAND2_X1 _1490_ (
  .A1(_0374_),
  .A2(_1234_),
  .ZN(_0383_)
);

INV_X1 _1491_ (
  .A(\ext_mult_res[7] ),
  .ZN(_0384_)
);

OAI21_X1 _1492_ (
  .A(_0383_),
  .B1(_0384_),
  .B2(_0372_),
  .ZN(_0007_)
);

INV_X1 _1493_ (
  .A(_0367_),
  .ZN(_0385_)
);

NAND2_X1 _1494_ (
  .A1(_0385_),
  .A2(\ext_mult_res[8] ),
  .ZN(_0386_)
);

BUF_X1 _1495_ (
  .A(_0385_),
  .Z(_0387_)
);

OAI21_X1 _1496_ (
  .A(_0386_),
  .B1(_0794_),
  .B2(_0387_),
  .ZN(_0008_)
);

INV_X1 _1497_ (
  .A(_0793_),
  .ZN(_0388_)
);

NAND2_X1 _1498_ (
  .A1(_0388_),
  .A2(_1185_),
  .ZN(_0389_)
);

INV_X1 _1499_ (
  .A(_1185_),
  .ZN(_0390_)
);

NAND2_X1 _1500_ (
  .A1(_0390_),
  .A2(_0793_),
  .ZN(_0391_)
);

NAND3_X1 _1501_ (
  .A1(_0389_),
  .A2(_0391_),
  .A3(_0374_),
  .ZN(_0392_)
);

INV_X1 _1502_ (
  .A(\ext_mult_res[9] ),
  .ZN(_0393_)
);

OAI21_X1 _1503_ (
  .A(_0392_),
  .B1(_0393_),
  .B2(_0372_),
  .ZN(_0009_)
);

NOR2_X1 _1504_ (
  .A1(\ext_mult_res[10] ),
  .A2(_0373_),
  .ZN(_0394_)
);

INV_X1 _1505_ (
  .A(_1184_),
  .ZN(_0395_)
);

INV_X1 _1506_ (
  .A(_1174_),
  .ZN(_0396_)
);

OAI21_X1 _1507_ (
  .A(_0395_),
  .B1(_0390_),
  .B2(_0396_),
  .ZN(_0397_)
);

INV_X1 _1508_ (
  .A(_0397_),
  .ZN(_0398_)
);

NAND2_X1 _1509_ (
  .A1(_1185_),
  .A2(_1175_),
  .ZN(_0399_)
);

OAI21_X1 _1510_ (
  .A(_0398_),
  .B1(_0792_),
  .B2(_0399_),
  .ZN(_0400_)
);

BUF_X1 _1511_ (
  .A(_1191_),
  .Z(_0401_)
);

XNOR2_X1 _1512_ (
  .A(_0400_),
  .B(_0401_),
  .ZN(_0402_)
);

BUF_X1 _1513_ (
  .A(_0371_),
  .Z(_0403_)
);

AOI21_X1 _1514_ (
  .A(_0394_),
  .B1(_0402_),
  .B2(_0403_),
  .ZN(_0010_)
);

NOR2_X1 _1515_ (
  .A1(\ext_mult_res[11] ),
  .A2(_0373_),
  .ZN(_0404_)
);

INV_X1 _1516_ (
  .A(_1190_),
  .ZN(_0405_)
);

INV_X1 _1517_ (
  .A(_0401_),
  .ZN(_0406_)
);

OAI21_X1 _1518_ (
  .A(_0405_),
  .B1(_0406_),
  .B2(_0395_),
  .ZN(_0407_)
);

NAND2_X1 _1519_ (
  .A1(_1185_),
  .A2(_0401_),
  .ZN(_0408_)
);

INV_X1 _1520_ (
  .A(_0408_),
  .ZN(_0409_)
);

AOI21_X1 _1521_ (
  .A(_0407_),
  .B1(_0409_),
  .B2(_0388_),
  .ZN(_0410_)
);

INV_X1 _1522_ (
  .A(_1198_),
  .ZN(_0411_)
);

XNOR2_X1 _1523_ (
  .A(_0410_),
  .B(_0411_),
  .ZN(_0412_)
);

AOI21_X1 _1524_ (
  .A(_0404_),
  .B1(_0412_),
  .B2(_0403_),
  .ZN(_0011_)
);

NOR2_X1 _1525_ (
  .A1(\ext_mult_res[12] ),
  .A2(_0373_),
  .ZN(_0413_)
);

INV_X1 _1526_ (
  .A(_1197_),
  .ZN(_0414_)
);

OAI21_X1 _1527_ (
  .A(_0414_),
  .B1(_0411_),
  .B2(_0405_),
  .ZN(_0415_)
);

INV_X1 _1528_ (
  .A(_0415_),
  .ZN(_0416_)
);

NAND2_X1 _1529_ (
  .A1(_0401_),
  .A2(_1198_),
  .ZN(_0417_)
);

OAI21_X1 _1530_ (
  .A(_0416_),
  .B1(_0398_),
  .B2(_0417_),
  .ZN(_0418_)
);

NOR2_X1 _1531_ (
  .A1(_0399_),
  .A2(_0417_),
  .ZN(_0419_)
);

AOI21_X1 _1532_ (
  .A(_0418_),
  .B1(_0419_),
  .B2(_1177_),
  .ZN(_0420_)
);

INV_X1 _1533_ (
  .A(_1203_),
  .ZN(_0421_)
);

XNOR2_X1 _1534_ (
  .A(_0420_),
  .B(_0421_),
  .ZN(_0422_)
);

AOI21_X1 _1535_ (
  .A(_0413_),
  .B1(_0422_),
  .B2(_0403_),
  .ZN(_0012_)
);

NOR2_X1 _1536_ (
  .A1(\ext_mult_res[13] ),
  .A2(_0373_),
  .ZN(_0423_)
);

INV_X1 _1537_ (
  .A(_1202_),
  .ZN(_0424_)
);

OAI21_X1 _1538_ (
  .A(_0424_),
  .B1(_0421_),
  .B2(_0414_),
  .ZN(_0425_)
);

INV_X1 _1539_ (
  .A(_0425_),
  .ZN(_0426_)
);

INV_X1 _1540_ (
  .A(_0407_),
  .ZN(_0427_)
);

NAND2_X1 _1541_ (
  .A1(_1198_),
  .A2(_1203_),
  .ZN(_0428_)
);

OAI21_X1 _1542_ (
  .A(_0426_),
  .B1(_0427_),
  .B2(_0428_),
  .ZN(_0429_)
);

NOR2_X1 _1543_ (
  .A1(_0408_),
  .A2(_0428_),
  .ZN(_0430_)
);

AOI21_X1 _1544_ (
  .A(_0429_),
  .B1(_0430_),
  .B2(_0388_),
  .ZN(_0431_)
);

INV_X1 _1545_ (
  .A(_1209_),
  .ZN(_0432_)
);

XNOR2_X1 _1546_ (
  .A(_0431_),
  .B(_0432_),
  .ZN(_0433_)
);

AOI21_X1 _1547_ (
  .A(_0423_),
  .B1(_0433_),
  .B2(_0403_),
  .ZN(_0013_)
);

NOR2_X1 _1548_ (
  .A1(\ext_mult_res[14] ),
  .A2(_0373_),
  .ZN(_0434_)
);

INV_X1 _1549_ (
  .A(_1208_),
  .ZN(_0435_)
);

OAI21_X1 _1550_ (
  .A(_0435_),
  .B1(_0432_),
  .B2(_0424_),
  .ZN(_0436_)
);

INV_X1 _1551_ (
  .A(_0436_),
  .ZN(_0437_)
);

NAND2_X1 _1552_ (
  .A1(_1203_),
  .A2(_1209_),
  .ZN(_0438_)
);

OAI21_X1 _1553_ (
  .A(_0437_),
  .B1(_0416_),
  .B2(_0438_),
  .ZN(_0439_)
);

NOR2_X1 _1554_ (
  .A1(_0417_),
  .A2(_0438_),
  .ZN(_0440_)
);

AOI21_X1 _1555_ (
  .A(_0439_),
  .B1(_0440_),
  .B2(_0400_),
  .ZN(_0441_)
);

INV_X1 _1556_ (
  .A(_1215_),
  .ZN(_0442_)
);

XNOR2_X1 _1557_ (
  .A(_0441_),
  .B(_0442_),
  .ZN(_0443_)
);

AOI21_X1 _1558_ (
  .A(_0434_),
  .B1(_0443_),
  .B2(_0403_),
  .ZN(_0014_)
);

NAND2_X1 _1559_ (
  .A1(_1209_),
  .A2(_1215_),
  .ZN(_0444_)
);

NOR3_X1 _1560_ (
  .A1(_0410_),
  .A2(_0428_),
  .A3(_0444_),
  .ZN(_0445_)
);

INV_X1 _1561_ (
  .A(_1214_),
  .ZN(_0446_)
);

OAI21_X1 _1562_ (
  .A(_0446_),
  .B1(_0442_),
  .B2(_0435_),
  .ZN(_0447_)
);

INV_X1 _1563_ (
  .A(_0447_),
  .ZN(_0448_)
);

OAI21_X1 _1564_ (
  .A(_0448_),
  .B1(_0426_),
  .B2(_0444_),
  .ZN(_0449_)
);

OR2_X1 _1565_ (
  .A1(_0445_),
  .A2(_0449_),
  .ZN(_0450_)
);

BUF_X1 _1566_ (
  .A(_1221_),
  .Z(_0451_)
);

OR2_X1 _1567_ (
  .A1(_0450_),
  .A2(_0451_),
  .ZN(_0452_)
);

NAND2_X1 _1568_ (
  .A1(_0450_),
  .A2(_0451_),
  .ZN(_0453_)
);

NAND3_X1 _1569_ (
  .A1(_0452_),
  .A2(_0374_),
  .A3(_0453_),
  .ZN(_0454_)
);

INV_X1 _1570_ (
  .A(\ext_mult_res[15] ),
  .ZN(_0455_)
);

OAI21_X1 _1571_ (
  .A(_0454_),
  .B1(_0455_),
  .B2(_0372_),
  .ZN(_0015_)
);

NOR2_X1 _1572_ (
  .A1(\ext_mult_res[16] ),
  .A2(_0373_),
  .ZN(_0456_)
);

INV_X1 _1573_ (
  .A(_1220_),
  .ZN(_0457_)
);

INV_X1 _1574_ (
  .A(_0451_),
  .ZN(_0458_)
);

OAI21_X1 _1575_ (
  .A(_0457_),
  .B1(_0458_),
  .B2(_0446_),
  .ZN(_0459_)
);

INV_X1 _1576_ (
  .A(_0459_),
  .ZN(_0460_)
);

NAND2_X1 _1577_ (
  .A1(_1215_),
  .A2(_0451_),
  .ZN(_0461_)
);

OAI21_X1 _1578_ (
  .A(_0460_),
  .B1(_0437_),
  .B2(_0461_),
  .ZN(_0462_)
);

NOR2_X1 _1579_ (
  .A1(_0438_),
  .A2(_0461_),
  .ZN(_0463_)
);

AOI21_X1 _1580_ (
  .A(_0462_),
  .B1(_0463_),
  .B2(_0418_),
  .ZN(_0464_)
);

NAND3_X1 _1581_ (
  .A1(_0419_),
  .A2(_0463_),
  .A3(_1177_),
  .ZN(_0465_)
);

NAND2_X1 _1582_ (
  .A1(_0464_),
  .A2(_0465_),
  .ZN(_0466_)
);

BUF_X1 _1583_ (
  .A(_1230_),
  .Z(_0467_)
);

XNOR2_X1 _1584_ (
  .A(_0466_),
  .B(_0467_),
  .ZN(_0468_)
);

AOI21_X1 _1585_ (
  .A(_0456_),
  .B1(_0468_),
  .B2(_0403_),
  .ZN(_0016_)
);

NOR2_X1 _1586_ (
  .A1(\ext_mult_res[17] ),
  .A2(_0373_),
  .ZN(_0469_)
);

INV_X1 _1587_ (
  .A(_1229_),
  .ZN(_0470_)
);

INV_X1 _1588_ (
  .A(_0467_),
  .ZN(_0471_)
);

NAND2_X1 _1589_ (
  .A1(_0451_),
  .A2(_0467_),
  .ZN(_0472_)
);

OAI221_X1 _1590_ (
  .A(_0470_),
  .B1(_0457_),
  .B2(_0471_),
  .C1(_0448_),
  .C2(_0472_),
  .ZN(_0473_)
);

INV_X1 _1591_ (
  .A(_0473_),
  .ZN(_0474_)
);

NOR2_X1 _1592_ (
  .A1(_0444_),
  .A2(_0472_),
  .ZN(_0475_)
);

NAND2_X1 _1593_ (
  .A1(_0429_),
  .A2(_0475_),
  .ZN(_0476_)
);

NAND3_X1 _1594_ (
  .A1(_0430_),
  .A2(_0475_),
  .A3(_0388_),
  .ZN(_0477_)
);

NAND3_X1 _1595_ (
  .A1(_0474_),
  .A2(_0476_),
  .A3(_0477_),
  .ZN(_0478_)
);

BUF_X1 _1596_ (
  .A(_1233_),
  .Z(_0479_)
);

XNOR2_X1 _1597_ (
  .A(_0478_),
  .B(_0479_),
  .ZN(_0480_)
);

AOI21_X1 _1598_ (
  .A(_0469_),
  .B1(_0480_),
  .B2(_0403_),
  .ZN(_0017_)
);

INV_X1 _1599_ (
  .A(_1061_),
  .ZN(_0481_)
);

INV_X1 _1600_ (
  .A(_1070_),
  .ZN(_0482_)
);

NAND2_X1 _1601_ (
  .A1(_0481_),
  .A2(_0482_),
  .ZN(_0483_)
);

NAND2_X1 _1602_ (
  .A1(_1061_),
  .A2(_1070_),
  .ZN(_0484_)
);

NAND2_X1 _1603_ (
  .A1(_0483_),
  .A2(_0484_),
  .ZN(_0485_)
);

INV_X1 _1604_ (
  .A(_0485_),
  .ZN(_0486_)
);

INV_X1 _1605_ (
  .A(_1081_),
  .ZN(_0487_)
);

NAND2_X1 _1606_ (
  .A1(_0487_),
  .A2(_1055_),
  .ZN(_0488_)
);

INV_X1 _1607_ (
  .A(_1055_),
  .ZN(_0489_)
);

NAND2_X1 _1608_ (
  .A1(_0489_),
  .A2(_1081_),
  .ZN(_0490_)
);

NAND2_X1 _1609_ (
  .A1(_0488_),
  .A2(_0490_),
  .ZN(_0491_)
);

NAND2_X1 _1610_ (
  .A1(_0486_),
  .A2(_0491_),
  .ZN(_0492_)
);

XNOR2_X1 _1611_ (
  .A(_1081_),
  .B(_1055_),
  .ZN(_0493_)
);

NAND2_X1 _1612_ (
  .A1(_0493_),
  .A2(_0485_),
  .ZN(_0494_)
);

NAND2_X1 _1613_ (
  .A1(_0492_),
  .A2(_0494_),
  .ZN(_0495_)
);

INV_X1 _1614_ (
  .A(_1224_),
  .ZN(_0496_)
);

NAND2_X1 _1615_ (
  .A1(_0496_),
  .A2(_1027_),
  .ZN(_0497_)
);

NAND2_X1 _1616_ (
  .A1(_1224_),
  .A2(_0987_),
  .ZN(_0498_)
);

NAND2_X1 _1617_ (
  .A1(_0497_),
  .A2(_0498_),
  .ZN(_0499_)
);

NAND2_X1 _1618_ (
  .A1(_0499_),
  .A2(_1023_),
  .ZN(_0500_)
);

NAND3_X1 _1619_ (
  .A1(_0497_),
  .A2(_1052_),
  .A3(_0498_),
  .ZN(_0501_)
);

NAND2_X2 _1620_ (
  .A1(_0500_),
  .A2(_0501_),
  .ZN(_0502_)
);

XNOR2_X1 _1621_ (
  .A(_0495_),
  .B(_0502_),
  .ZN(_0503_)
);

INV_X1 _1622_ (
  .A(_1005_),
  .ZN(_0504_)
);

XNOR2_X1 _1623_ (
  .A(_0504_),
  .B(_1059_),
  .ZN(_0505_)
);

XNOR2_X1 _1624_ (
  .A(_1063_),
  .B(_1065_),
  .ZN(_0506_)
);

NAND2_X1 _1625_ (
  .A1(_0505_),
  .A2(_0506_),
  .ZN(_0507_)
);

NAND2_X1 _1626_ (
  .A1(_1063_),
  .A2(_1065_),
  .ZN(_0508_)
);

INV_X1 _1627_ (
  .A(_0508_),
  .ZN(_0509_)
);

NOR2_X1 _1628_ (
  .A1(_1063_),
  .A2(_1065_),
  .ZN(_0510_)
);

NOR2_X1 _1629_ (
  .A1(_0509_),
  .A2(_0510_),
  .ZN(_0511_)
);

XNOR2_X1 _1630_ (
  .A(_1005_),
  .B(_1059_),
  .ZN(_0512_)
);

NAND2_X1 _1631_ (
  .A1(_0511_),
  .A2(_0512_),
  .ZN(_0513_)
);

NAND2_X1 _1632_ (
  .A1(_0507_),
  .A2(_0513_),
  .ZN(_0514_)
);

INV_X1 _1633_ (
  .A(_0514_),
  .ZN(_0515_)
);

NAND2_X2 _1637_ (
  .A1(_0518_),
  .A2(_1053_),
  .ZN(_0519_)
);

NAND2_X2 _1639_ (
  .A1(_0519_),
  .A2(_0520_),
  .ZN(_0521_)
);

NAND2_X1 _1640_ (
  .A1(_0515_),
  .A2(_0521_),
  .ZN(_0522_)
);

NAND2_X2 _1641_ (
  .A1(_0518_),
  .A2(_1024_),
  .ZN(_0523_)
);

INV_X1 _1642_ (
  .A(_0358_),
  .ZN(_0524_)
);

NAND2_X2 _1644_ (
  .A1(_0523_),
  .A2(_0525_),
  .ZN(_0526_)
);

NAND2_X1 _1645_ (
  .A1(_0526_),
  .A2(_0514_),
  .ZN(_0527_)
);

NAND2_X2 _1646_ (
  .A1(_0522_),
  .A2(_0527_),
  .ZN(_0528_)
);

NAND2_X1 _1647_ (
  .A1(_0503_),
  .A2(_0528_),
  .ZN(_0529_)
);

NAND2_X1 _1648_ (
  .A1(_0515_),
  .A2(_0526_),
  .ZN(_0530_)
);

NAND2_X1 _1649_ (
  .A1(_0521_),
  .A2(_0514_),
  .ZN(_0531_)
);

NAND2_X2 _1650_ (
  .A1(_0530_),
  .A2(_0531_),
  .ZN(_0532_)
);

XNOR2_X1 _1651_ (
  .A(_0491_),
  .B(_0485_),
  .ZN(_0533_)
);

NAND2_X1 _1652_ (
  .A1(_0533_),
  .A2(_0502_),
  .ZN(_0534_)
);

INV_X1 _1653_ (
  .A(_0502_),
  .ZN(_0535_)
);

NAND2_X1 _1654_ (
  .A1(_0495_),
  .A2(_0535_),
  .ZN(_0536_)
);

NAND2_X1 _1655_ (
  .A1(_0534_),
  .A2(_0536_),
  .ZN(_0537_)
);

NAND2_X1 _1656_ (
  .A1(_0532_),
  .A2(_0537_),
  .ZN(_0538_)
);

NAND2_X1 _1657_ (
  .A1(_0529_),
  .A2(_0538_),
  .ZN(_0539_)
);

OR2_X1 _1658_ (
  .A1(_1086_),
  .A2(_1078_),
  .ZN(_0540_)
);

NAND2_X1 _1659_ (
  .A1(_1078_),
  .A2(_1086_),
  .ZN(_0541_)
);

XOR2_X1 _1664_ (
  .A(_1068_),
  .B(_1231_),
  .Z(_0546_)
);

INV_X1 _1665_ (
  .A(_0546_),
  .ZN(_0547_)
);

NAND2_X2 _1666_ (
  .A1(_0545_),
  .A2(_0547_),
  .ZN(_0548_)
);

NAND2_X2 _1668_ (
  .A1(_0548_),
  .A2(_0549_),
  .ZN(_0550_)
);

XNOR2_X1 _1669_ (
  .A(_0967_),
  .B(_0903_),
  .ZN(_0551_)
);

XNOR2_X1 _1670_ (
  .A(_0874_),
  .B(_1073_),
  .ZN(_0552_)
);

XNOR2_X1 _1671_ (
  .A(_0551_),
  .B(_0552_),
  .ZN(_0553_)
);

INV_X1 _1672_ (
  .A(_0553_),
  .ZN(_0554_)
);

NAND2_X2 _1673_ (
  .A1(_0550_),
  .A2(_0554_),
  .ZN(_0555_)
);

NAND3_X1 _1674_ (
  .A1(_0548_),
  .A2(_0549_),
  .A3(_0553_),
  .ZN(_0556_)
);

NAND2_X2 _1675_ (
  .A1(_0555_),
  .A2(_0556_),
  .ZN(_0557_)
);

INV_X1 _1676_ (
  .A(_0557_),
  .ZN(_0558_)
);

NAND2_X2 _1677_ (
  .A1(_0539_),
  .A2(_0558_),
  .ZN(_0559_)
);

NAND2_X1 _1678_ (
  .A1(_0503_),
  .A2(_0532_),
  .ZN(_0560_)
);

NAND2_X1 _1679_ (
  .A1(_0528_),
  .A2(_0537_),
  .ZN(_0561_)
);

NAND2_X2 _1680_ (
  .A1(_0560_),
  .A2(_0561_),
  .ZN(_0562_)
);

NAND2_X2 _1681_ (
  .A1(_0562_),
  .A2(_0557_),
  .ZN(_0563_)
);

NAND2_X2 _1682_ (
  .A1(_0559_),
  .A2(_0563_),
  .ZN(_0564_)
);

INV_X1 _1683_ (
  .A(_0479_),
  .ZN(_0565_)
);

NOR3_X1 _1684_ (
  .A1(_0461_),
  .A2(_0471_),
  .A3(_0565_),
  .ZN(_0566_)
);

NAND3_X1 _1685_ (
  .A1(_0400_),
  .A2(_0440_),
  .A3(_0566_),
  .ZN(_0567_)
);

NAND3_X1 _1686_ (
  .A1(_0459_),
  .A2(_0467_),
  .A3(_0479_),
  .ZN(_0568_)
);

INV_X1 _1687_ (
  .A(_1232_),
  .ZN(_0569_)
);

NAND2_X1 _1688_ (
  .A1(_0479_),
  .A2(_1229_),
  .ZN(_0570_)
);

NAND3_X1 _1689_ (
  .A1(_0568_),
  .A2(_0569_),
  .A3(_0570_),
  .ZN(_0571_)
);

INV_X1 _1690_ (
  .A(_0571_),
  .ZN(_0572_)
);

NAND2_X1 _1691_ (
  .A1(_0439_),
  .A2(_0566_),
  .ZN(_0573_)
);

AND3_X1 _1692_ (
  .A1(_0567_),
  .A2(_0572_),
  .A3(_0573_),
  .ZN(_0574_)
);

INV_X1 _1693_ (
  .A(_0574_),
  .ZN(_0575_)
);

NAND2_X2 _1694_ (
  .A1(_0564_),
  .A2(_0575_),
  .ZN(_0576_)
);

NAND3_X1 _1695_ (
  .A1(_0559_),
  .A2(_0563_),
  .A3(_0574_),
  .ZN(_0577_)
);

NAND3_X1 _1696_ (
  .A1(_0576_),
  .A2(_0577_),
  .A3(_0374_),
  .ZN(_0578_)
);

NAND2_X1 _1697_ (
  .A1(_0387_),
  .A2(\ext_mult_res[18] ),
  .ZN(_0579_)
);

NAND2_X1 _1698_ (
  .A1(_0578_),
  .A2(_0579_),
  .ZN(_0018_)
);

NAND2_X1 _1699_ (
  .A1(_0385_),
  .A2(result[0]),
  .ZN(_0580_)
);

BUF_X1 _1700_ (
  .A(dclr),
  .Z(_0581_)
);

OAI21_X1 _1701_ (
  .A(_0368_),
  .B1(_1089_),
  .B2(_0581_),
  .ZN(_0582_)
);

INV_X1 _1702_ (
  .A(_0581_),
  .ZN(_0583_)
);

BUF_X1 _1703_ (
  .A(_0583_),
  .Z(_0584_)
);

NOR2_X1 _1704_ (
  .A1(_0584_),
  .A2(\ext_mult_res[0] ),
  .ZN(_0585_)
);

OAI21_X1 _1705_ (
  .A(_0580_),
  .B1(_0582_),
  .B2(_0585_),
  .ZN(_0019_)
);

NAND2_X1 _1706_ (
  .A1(_0385_),
  .A2(result[1]),
  .ZN(_0586_)
);

OAI21_X1 _1707_ (
  .A(_0368_),
  .B1(_0581_),
  .B2(_0680_),
  .ZN(_0587_)
);

NOR2_X1 _1708_ (
  .A1(_0584_),
  .A2(\ext_mult_res[1] ),
  .ZN(_0588_)
);

OAI21_X1 _1709_ (
  .A(_0586_),
  .B1(_0587_),
  .B2(_0588_),
  .ZN(_0020_)
);

INV_X1 _1710_ (
  .A(_1093_),
  .ZN(_0589_)
);

NOR2_X1 _1711_ (
  .A1(_0589_),
  .A2(_0679_),
  .ZN(_0590_)
);

INV_X1 _1712_ (
  .A(_0590_),
  .ZN(_0591_)
);

NAND2_X1 _1713_ (
  .A1(_0589_),
  .A2(_0679_),
  .ZN(_0592_)
);

NAND3_X1 _1714_ (
  .A1(_0591_),
  .A2(_0583_),
  .A3(_0592_),
  .ZN(_0593_)
);

BUF_X2 _1715_ (
  .A(_0583_),
  .Z(_0594_)
);

OAI21_X1 _1716_ (
  .A(_0593_),
  .B1(_0594_),
  .B2(_0376_),
  .ZN(_0595_)
);

MUX2_X1 _1717_ (
  .A(result[2]),
  .B(_0595_),
  .S(_0373_),
  .Z(_0021_)
);

OAI21_X1 _1718_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(_0378_),
  .ZN(_0596_)
);

NAND2_X1 _1719_ (
  .A1(_1088_),
  .A2(_1091_),
  .ZN(_0597_)
);

INV_X1 _1720_ (
  .A(_1090_),
  .ZN(_0598_)
);

INV_X1 _1721_ (
  .A(_1092_),
  .ZN(_0599_)
);

NAND3_X1 _1722_ (
  .A1(_0597_),
  .A2(_0598_),
  .A3(_0599_),
  .ZN(_0600_)
);

NAND2_X1 _1723_ (
  .A1(_0589_),
  .A2(_0599_),
  .ZN(_0601_)
);

NAND2_X1 _1724_ (
  .A1(_0600_),
  .A2(_0601_),
  .ZN(_0602_)
);

XNOR2_X1 _1725_ (
  .A(_0602_),
  .B(_1095_),
  .ZN(_0603_)
);

BUF_X1 _1726_ (
  .A(_0583_),
  .Z(_0604_)
);

AOI21_X1 _1727_ (
  .A(_0596_),
  .B1(_0603_),
  .B2(_0604_),
  .ZN(_0605_)
);

INV_X1 _1728_ (
  .A(result[3]),
  .ZN(_0606_)
);

AOI21_X1 _1729_ (
  .A(_0605_),
  .B1(_0606_),
  .B2(_0387_),
  .ZN(_0022_)
);

OAI21_X1 _1730_ (
  .A(_0367_),
  .B1(_0583_),
  .B2(_0380_),
  .ZN(_0607_)
);

INV_X1 _1731_ (
  .A(_1094_),
  .ZN(_0608_)
);

INV_X1 _1732_ (
  .A(_1095_),
  .ZN(_0609_)
);

OAI21_X1 _1733_ (
  .A(_0608_),
  .B1(_0609_),
  .B2(_0599_),
  .ZN(_0610_)
);

INV_X1 _1734_ (
  .A(_0610_),
  .ZN(_0611_)
);

OAI21_X4 _1735_ (
  .A(_0611_),
  .B1(_0609_),
  .B2(_0591_),
  .ZN(_0612_)
);

INV_X1 _1736_ (
  .A(_1097_),
  .ZN(_0613_)
);

XNOR2_X1 _1737_ (
  .A(_0612_),
  .B(_0613_),
  .ZN(_0614_)
);

AOI21_X1 _1738_ (
  .A(_0607_),
  .B1(_0614_),
  .B2(_0604_),
  .ZN(_0615_)
);

INV_X1 _1739_ (
  .A(result[4]),
  .ZN(_0616_)
);

AOI21_X1 _1740_ (
  .A(_0615_),
  .B1(_0616_),
  .B2(_0387_),
  .ZN(_0023_)
);

NAND2_X1 _1741_ (
  .A1(_1095_),
  .A2(_1097_),
  .ZN(_0617_)
);

INV_X1 _1742_ (
  .A(_0617_),
  .ZN(_0618_)
);

NAND3_X1 _1743_ (
  .A1(_0600_),
  .A2(_0601_),
  .A3(_0618_),
  .ZN(_0619_)
);

INV_X1 _1744_ (
  .A(_1096_),
  .ZN(_0620_)
);

OAI21_X1 _1745_ (
  .A(_0620_),
  .B1(_0613_),
  .B2(_0608_),
  .ZN(_0621_)
);

INV_X1 _1746_ (
  .A(_0621_),
  .ZN(_0622_)
);

NAND2_X1 _1747_ (
  .A1(_0619_),
  .A2(_0622_),
  .ZN(_0623_)
);

BUF_X2 _1748_ (
  .A(_1099_),
  .Z(_0624_)
);

XNOR2_X1 _1749_ (
  .A(_0623_),
  .B(_0624_),
  .ZN(_0625_)
);

AOI21_X1 _1750_ (
  .A(_0385_),
  .B1(_0625_),
  .B2(_0594_),
  .ZN(_0626_)
);

OAI21_X1 _1751_ (
  .A(_0626_),
  .B1(_0584_),
  .B2(\ext_mult_res[5] ),
  .ZN(_0627_)
);

INV_X1 _1752_ (
  .A(result[5]),
  .ZN(_0628_)
);

OAI21_X1 _1753_ (
  .A(_0627_),
  .B1(_0403_),
  .B2(_0628_),
  .ZN(_0024_)
);

INV_X1 _1754_ (
  .A(_1098_),
  .ZN(_0629_)
);

INV_X1 _1755_ (
  .A(_0624_),
  .ZN(_0630_)
);

OAI21_X1 _1756_ (
  .A(_0629_),
  .B1(_0630_),
  .B2(_0620_),
  .ZN(_0631_)
);

INV_X1 _1757_ (
  .A(_0631_),
  .ZN(_0632_)
);

INV_X1 _1758_ (
  .A(_0612_),
  .ZN(_0633_)
);

NAND2_X1 _1759_ (
  .A1(_1097_),
  .A2(_0624_),
  .ZN(_0634_)
);

OAI21_X1 _1760_ (
  .A(_0632_),
  .B1(_0633_),
  .B2(_0634_),
  .ZN(_0635_)
);

CLKBUF_X2 _1761_ (
  .A(_1101_),
  .Z(_0636_)
);

XNOR2_X1 _1762_ (
  .A(_0635_),
  .B(_0636_),
  .ZN(_0041_)
);

NAND2_X1 _1763_ (
  .A1(_0041_),
  .A2(_0604_),
  .ZN(_0042_)
);

NAND2_X1 _1764_ (
  .A1(_0382_),
  .A2(_0581_),
  .ZN(_0043_)
);

NAND3_X1 _1765_ (
  .A1(_0042_),
  .A2(_0374_),
  .A3(_0043_),
  .ZN(_0044_)
);

INV_X1 _1766_ (
  .A(result[6]),
  .ZN(_0045_)
);

OAI21_X1 _1767_ (
  .A(_0044_),
  .B1(_0403_),
  .B2(_0045_),
  .ZN(_0025_)
);

NAND2_X1 _1768_ (
  .A1(_0636_),
  .A2(_1098_),
  .ZN(_0046_)
);

INV_X1 _1769_ (
  .A(_1100_),
  .ZN(_0047_)
);

NAND2_X1 _1770_ (
  .A1(_0046_),
  .A2(_0047_),
  .ZN(_0048_)
);

INV_X1 _1771_ (
  .A(_0048_),
  .ZN(_0049_)
);

NAND2_X1 _1772_ (
  .A1(_0624_),
  .A2(_0636_),
  .ZN(_0050_)
);

OAI21_X1 _1773_ (
  .A(_0049_),
  .B1(_0622_),
  .B2(_0050_),
  .ZN(_0051_)
);

INV_X1 _1774_ (
  .A(_0051_),
  .ZN(_0052_)
);

OAI21_X1 _1775_ (
  .A(_0052_),
  .B1(_0619_),
  .B2(_0050_),
  .ZN(_0053_)
);

BUF_X2 _1776_ (
  .A(_1103_),
  .Z(_0054_)
);

XNOR2_X1 _1777_ (
  .A(_0053_),
  .B(_0054_),
  .ZN(_0055_)
);

NAND2_X1 _1778_ (
  .A1(_0055_),
  .A2(_0604_),
  .ZN(_0056_)
);

NAND2_X1 _1779_ (
  .A1(_0384_),
  .A2(_0581_),
  .ZN(_0057_)
);

NAND3_X1 _1780_ (
  .A1(_0056_),
  .A2(_0374_),
  .A3(_0057_),
  .ZN(_0058_)
);

INV_X1 _1781_ (
  .A(result[7]),
  .ZN(_0059_)
);

OAI21_X1 _1782_ (
  .A(_0058_),
  .B1(_0403_),
  .B2(_0059_),
  .ZN(_0026_)
);

NAND2_X1 _1783_ (
  .A1(_0385_),
  .A2(result[8]),
  .ZN(_0060_)
);

INV_X1 _1784_ (
  .A(_1102_),
  .ZN(_0061_)
);

INV_X1 _1785_ (
  .A(_0054_),
  .ZN(_0062_)
);

OAI21_X1 _1786_ (
  .A(_0061_),
  .B1(_0062_),
  .B2(_0047_),
  .ZN(_0063_)
);

INV_X1 _1787_ (
  .A(_0063_),
  .ZN(_0064_)
);

NAND2_X1 _1788_ (
  .A1(_0636_),
  .A2(_0054_),
  .ZN(_0065_)
);

OAI21_X1 _1789_ (
  .A(_0064_),
  .B1(_0632_),
  .B2(_0065_),
  .ZN(_0066_)
);

INV_X1 _1790_ (
  .A(_0066_),
  .ZN(_0067_)
);

NOR2_X1 _1791_ (
  .A1(_0634_),
  .A2(_0065_),
  .ZN(_0068_)
);

INV_X1 _1792_ (
  .A(_0068_),
  .ZN(_0069_)
);

OAI21_X1 _1793_ (
  .A(_0067_),
  .B1(_0633_),
  .B2(_0069_),
  .ZN(_0070_)
);

INV_X1 _1794_ (
  .A(_1105_),
  .ZN(_0071_)
);

XNOR2_X1 _1795_ (
  .A(_0070_),
  .B(_0071_),
  .ZN(_0072_)
);

OAI21_X1 _1796_ (
  .A(_0368_),
  .B1(_0072_),
  .B2(_0581_),
  .ZN(_0073_)
);

NOR2_X1 _1797_ (
  .A1(_0584_),
  .A2(\ext_mult_res[8] ),
  .ZN(_0074_)
);

OAI21_X1 _1798_ (
  .A(_0060_),
  .B1(_0073_),
  .B2(_0074_),
  .ZN(_0027_)
);

OAI21_X1 _1799_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[9] ),
  .ZN(_0075_)
);

INV_X1 _1800_ (
  .A(_0075_),
  .ZN(_0076_)
);

NAND2_X2 _1801_ (
  .A1(_0054_),
  .A2(_1105_),
  .ZN(_0077_)
);

INV_X1 _1802_ (
  .A(_0077_),
  .ZN(_0078_)
);

NAND2_X1 _1803_ (
  .A1(_0053_),
  .A2(_0078_),
  .ZN(_0079_)
);

INV_X1 _1804_ (
  .A(_1104_),
  .ZN(_0080_)
);

OAI21_X1 _1805_ (
  .A(_0080_),
  .B1(_0071_),
  .B2(_0061_),
  .ZN(_0081_)
);

INV_X1 _1806_ (
  .A(_0081_),
  .ZN(_0082_)
);

NAND2_X1 _1807_ (
  .A1(_0079_),
  .A2(_0082_),
  .ZN(_0083_)
);

INV_X1 _1808_ (
  .A(_1107_),
  .ZN(_0084_)
);

XNOR2_X1 _1809_ (
  .A(_0083_),
  .B(_0084_),
  .ZN(_0085_)
);

OAI21_X1 _1810_ (
  .A(_0076_),
  .B1(_0085_),
  .B2(_0581_),
  .ZN(_0086_)
);

NAND2_X1 _1811_ (
  .A1(_0387_),
  .A2(result[9]),
  .ZN(_0087_)
);

NAND2_X1 _1812_ (
  .A1(_0086_),
  .A2(_0087_),
  .ZN(_0028_)
);

NAND2_X1 _1813_ (
  .A1(_0385_),
  .A2(result[10]),
  .ZN(_0088_)
);

OAI21_X1 _1814_ (
  .A(_0632_),
  .B1(_0611_),
  .B2(_0634_),
  .ZN(_0089_)
);

NAND2_X1 _1815_ (
  .A1(_1105_),
  .A2(_1107_),
  .ZN(_0090_)
);

NOR2_X1 _1816_ (
  .A1(_0065_),
  .A2(_0090_),
  .ZN(_0091_)
);

NAND2_X1 _1817_ (
  .A1(_0089_),
  .A2(_0091_),
  .ZN(_0092_)
);

INV_X1 _1818_ (
  .A(_1106_),
  .ZN(_0093_)
);

OAI21_X1 _1819_ (
  .A(_0093_),
  .B1(_0084_),
  .B2(_0080_),
  .ZN(_0094_)
);

INV_X1 _1820_ (
  .A(_0094_),
  .ZN(_0095_)
);

OAI21_X1 _1821_ (
  .A(_0095_),
  .B1(_0064_),
  .B2(_0090_),
  .ZN(_0096_)
);

INV_X1 _1822_ (
  .A(_0096_),
  .ZN(_0097_)
);

NOR3_X1 _1823_ (
  .A1(_0634_),
  .A2(_0589_),
  .A3(_0609_),
  .ZN(_0098_)
);

INV_X1 _1824_ (
  .A(_0679_),
  .ZN(_0099_)
);

NAND3_X1 _1825_ (
  .A1(_0098_),
  .A2(_0099_),
  .A3(_0091_),
  .ZN(_0100_)
);

NAND3_X1 _1826_ (
  .A1(_0092_),
  .A2(_0097_),
  .A3(_0100_),
  .ZN(_0101_)
);

INV_X1 _1827_ (
  .A(_1109_),
  .ZN(_0102_)
);

XNOR2_X1 _1828_ (
  .A(_0101_),
  .B(_0102_),
  .ZN(_0103_)
);

NOR2_X1 _1829_ (
  .A1(_0103_),
  .A2(_0581_),
  .ZN(_0104_)
);

OAI21_X1 _1830_ (
  .A(_0368_),
  .B1(_0584_),
  .B2(\ext_mult_res[10] ),
  .ZN(_0105_)
);

OAI21_X1 _1831_ (
  .A(_0088_),
  .B1(_0104_),
  .B2(_0105_),
  .ZN(_0029_)
);

NAND2_X1 _1832_ (
  .A1(_0385_),
  .A2(result[11]),
  .ZN(_0106_)
);

NAND2_X1 _1833_ (
  .A1(_1107_),
  .A2(_1109_),
  .ZN(_0107_)
);

NOR2_X2 _1834_ (
  .A1(_0077_),
  .A2(_0107_),
  .ZN(_0108_)
);

NAND2_X1 _1835_ (
  .A1(_0051_),
  .A2(_0108_),
  .ZN(_0109_)
);

INV_X1 _1836_ (
  .A(_1108_),
  .ZN(_0110_)
);

OAI21_X1 _1837_ (
  .A(_0110_),
  .B1(_0102_),
  .B2(_0093_),
  .ZN(_0111_)
);

INV_X1 _1838_ (
  .A(_0111_),
  .ZN(_0112_)
);

OAI21_X1 _1839_ (
  .A(_0112_),
  .B1(_0082_),
  .B2(_0107_),
  .ZN(_0113_)
);

INV_X1 _1840_ (
  .A(_0113_),
  .ZN(_0114_)
);

NAND2_X1 _1841_ (
  .A1(_0109_),
  .A2(_0114_),
  .ZN(_0115_)
);

INV_X1 _1842_ (
  .A(_0115_),
  .ZN(_0116_)
);

NAND4_X1 _1843_ (
  .A1(_0108_),
  .A2(_0618_),
  .A3(_0636_),
  .A4(_0624_),
  .ZN(_0117_)
);

INV_X1 _1844_ (
  .A(_0117_),
  .ZN(_0118_)
);

INV_X1 _1845_ (
  .A(_0602_),
  .ZN(_0119_)
);

NAND2_X1 _1846_ (
  .A1(_0118_),
  .A2(_0119_),
  .ZN(_0120_)
);

NAND2_X1 _1847_ (
  .A1(_0116_),
  .A2(_0120_),
  .ZN(_0121_)
);

INV_X1 _1848_ (
  .A(_1111_),
  .ZN(_0122_)
);

NAND2_X1 _1849_ (
  .A1(_0121_),
  .A2(_0122_),
  .ZN(_0123_)
);

NAND3_X1 _1850_ (
  .A1(_0116_),
  .A2(_1111_),
  .A3(_0120_),
  .ZN(_0124_)
);

NAND3_X1 _1851_ (
  .A1(_0123_),
  .A2(_0124_),
  .A3(_0604_),
  .ZN(_0125_)
);

NAND2_X1 _1852_ (
  .A1(_0125_),
  .A2(_0374_),
  .ZN(_0126_)
);

NOR2_X1 _1853_ (
  .A1(_0584_),
  .A2(\ext_mult_res[11] ),
  .ZN(_0127_)
);

OAI21_X1 _1854_ (
  .A(_0106_),
  .B1(_0126_),
  .B2(_0127_),
  .ZN(_0030_)
);

NAND2_X1 _1855_ (
  .A1(_0385_),
  .A2(result[12]),
  .ZN(_0128_)
);

NAND2_X1 _1856_ (
  .A1(_1109_),
  .A2(_1111_),
  .ZN(_0129_)
);

NOR2_X1 _1857_ (
  .A1(_0090_),
  .A2(_0129_),
  .ZN(_0130_)
);

NAND2_X1 _1858_ (
  .A1(_0066_),
  .A2(_0130_),
  .ZN(_0131_)
);

INV_X1 _1859_ (
  .A(_1110_),
  .ZN(_0132_)
);

OAI21_X1 _1860_ (
  .A(_0132_),
  .B1(_0122_),
  .B2(_0110_),
  .ZN(_0133_)
);

INV_X1 _1861_ (
  .A(_0133_),
  .ZN(_0134_)
);

OAI21_X1 _1862_ (
  .A(_0134_),
  .B1(_0095_),
  .B2(_0129_),
  .ZN(_0135_)
);

INV_X1 _1863_ (
  .A(_0135_),
  .ZN(_0136_)
);

NAND2_X1 _1864_ (
  .A1(_0131_),
  .A2(_0136_),
  .ZN(_0137_)
);

INV_X1 _1865_ (
  .A(_0137_),
  .ZN(_0138_)
);

NAND2_X1 _1866_ (
  .A1(_0068_),
  .A2(_0130_),
  .ZN(_0139_)
);

INV_X1 _1867_ (
  .A(_0139_),
  .ZN(_0140_)
);

NAND2_X1 _1868_ (
  .A1(_0612_),
  .A2(_0140_),
  .ZN(_0141_)
);

NAND2_X1 _1869_ (
  .A1(_0138_),
  .A2(_0141_),
  .ZN(_0142_)
);

INV_X1 _1870_ (
  .A(_1113_),
  .ZN(_0143_)
);

NAND2_X1 _1871_ (
  .A1(_0142_),
  .A2(_0143_),
  .ZN(_0144_)
);

NAND3_X1 _1872_ (
  .A1(_0138_),
  .A2(_1113_),
  .A3(_0141_),
  .ZN(_0145_)
);

AND3_X1 _1873_ (
  .A1(_0144_),
  .A2(_0145_),
  .A3(_0594_),
  .ZN(_0146_)
);

OAI21_X1 _1874_ (
  .A(_0368_),
  .B1(_0584_),
  .B2(\ext_mult_res[12] ),
  .ZN(_0147_)
);

OAI21_X1 _1875_ (
  .A(_0128_),
  .B1(_0146_),
  .B2(_0147_),
  .ZN(_0031_)
);

NAND2_X1 _1876_ (
  .A1(_0385_),
  .A2(result[13]),
  .ZN(_0148_)
);

NAND2_X1 _1877_ (
  .A1(_0048_),
  .A2(_0078_),
  .ZN(_0149_)
);

NAND2_X1 _1878_ (
  .A1(_0082_),
  .A2(_0149_),
  .ZN(_0150_)
);

NAND2_X1 _1879_ (
  .A1(_1111_),
  .A2(_1113_),
  .ZN(_0151_)
);

NOR2_X1 _1880_ (
  .A1(_0107_),
  .A2(_0151_),
  .ZN(_0152_)
);

NAND2_X1 _1881_ (
  .A1(_0150_),
  .A2(_0152_),
  .ZN(_0153_)
);

INV_X1 _1882_ (
  .A(_0151_),
  .ZN(_0154_)
);

NAND2_X1 _1883_ (
  .A1(_0111_),
  .A2(_0154_),
  .ZN(_0155_)
);

INV_X1 _1884_ (
  .A(_1112_),
  .ZN(_0156_)
);

OAI21_X1 _1885_ (
  .A(_0156_),
  .B1(_0143_),
  .B2(_0132_),
  .ZN(_0157_)
);

INV_X1 _1886_ (
  .A(_0157_),
  .ZN(_0158_)
);

NAND2_X1 _1887_ (
  .A1(_0155_),
  .A2(_0158_),
  .ZN(_0159_)
);

INV_X1 _1888_ (
  .A(_0159_),
  .ZN(_0160_)
);

NAND2_X1 _1889_ (
  .A1(_0153_),
  .A2(_0160_),
  .ZN(_0161_)
);

INV_X1 _1890_ (
  .A(_0161_),
  .ZN(_0162_)
);

INV_X1 _1891_ (
  .A(_0623_),
  .ZN(_0163_)
);

NOR2_X2 _1892_ (
  .A1(_0050_),
  .A2(_0077_),
  .ZN(_0164_)
);

NAND2_X1 _1893_ (
  .A1(_0164_),
  .A2(_0152_),
  .ZN(_0165_)
);

OAI21_X1 _1894_ (
  .A(_0162_),
  .B1(_0163_),
  .B2(_0165_),
  .ZN(_0166_)
);

INV_X1 _1895_ (
  .A(_1115_),
  .ZN(_0167_)
);

XNOR2_X1 _1896_ (
  .A(_0166_),
  .B(_0167_),
  .ZN(_0168_)
);

NOR2_X1 _1897_ (
  .A1(_0168_),
  .A2(_0581_),
  .ZN(_0169_)
);

OAI21_X1 _1898_ (
  .A(_0368_),
  .B1(_0604_),
  .B2(\ext_mult_res[13] ),
  .ZN(_0170_)
);

OAI21_X1 _1899_ (
  .A(_0148_),
  .B1(_0169_),
  .B2(_0170_),
  .ZN(_0032_)
);

NAND2_X1 _1900_ (
  .A1(_1113_),
  .A2(_1115_),
  .ZN(_0171_)
);

NOR2_X1 _1901_ (
  .A1(_0129_),
  .A2(_0171_),
  .ZN(_0172_)
);

NAND3_X1 _1902_ (
  .A1(_0635_),
  .A2(_0091_),
  .A3(_0172_),
  .ZN(_0173_)
);

INV_X1 _1903_ (
  .A(_1114_),
  .ZN(_0174_)
);

OAI21_X1 _1904_ (
  .A(_0174_),
  .B1(_0167_),
  .B2(_0156_),
  .ZN(_0175_)
);

INV_X1 _1905_ (
  .A(_0175_),
  .ZN(_0176_)
);

OAI21_X1 _1906_ (
  .A(_0176_),
  .B1(_0134_),
  .B2(_0171_),
  .ZN(_0177_)
);

AOI21_X1 _1907_ (
  .A(_0177_),
  .B1(_0172_),
  .B2(_0096_),
  .ZN(_0178_)
);

NAND2_X1 _1908_ (
  .A1(_0173_),
  .A2(_0178_),
  .ZN(_0179_)
);

INV_X1 _1909_ (
  .A(_1117_),
  .ZN(_0180_)
);

NAND2_X1 _1910_ (
  .A1(_0179_),
  .A2(_0180_),
  .ZN(_0181_)
);

NAND3_X1 _1911_ (
  .A1(_0173_),
  .A2(_1117_),
  .A3(_0178_),
  .ZN(_0182_)
);

NAND3_X1 _1912_ (
  .A1(_0181_),
  .A2(_0182_),
  .A3(_0604_),
  .ZN(_0183_)
);

OAI21_X1 _1913_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[14] ),
  .ZN(_0184_)
);

INV_X1 _1914_ (
  .A(_0184_),
  .ZN(_0185_)
);

NAND2_X1 _1915_ (
  .A1(_0183_),
  .A2(_0185_),
  .ZN(_0186_)
);

NAND2_X1 _1916_ (
  .A1(_0387_),
  .A2(result[14]),
  .ZN(_0187_)
);

NAND2_X1 _1917_ (
  .A1(_0186_),
  .A2(_0187_),
  .ZN(_0033_)
);

NAND2_X1 _1918_ (
  .A1(_1115_),
  .A2(_1117_),
  .ZN(_0188_)
);

NOR2_X1 _1919_ (
  .A1(_0151_),
  .A2(_0188_),
  .ZN(_0189_)
);

NAND3_X1 _1920_ (
  .A1(_0053_),
  .A2(_0108_),
  .A3(_0189_),
  .ZN(_0190_)
);

INV_X1 _1921_ (
  .A(_1116_),
  .ZN(_0191_)
);

OAI21_X1 _1922_ (
  .A(_0191_),
  .B1(_0180_),
  .B2(_0174_),
  .ZN(_0192_)
);

INV_X1 _1923_ (
  .A(_0192_),
  .ZN(_0193_)
);

OAI21_X1 _1924_ (
  .A(_0193_),
  .B1(_0158_),
  .B2(_0188_),
  .ZN(_0194_)
);

AOI21_X1 _1925_ (
  .A(_0194_),
  .B1(_0189_),
  .B2(_0113_),
  .ZN(_0195_)
);

NAND2_X1 _1926_ (
  .A1(_0190_),
  .A2(_0195_),
  .ZN(_0196_)
);

INV_X1 _1927_ (
  .A(_1119_),
  .ZN(_0197_)
);

NAND2_X1 _1928_ (
  .A1(_0196_),
  .A2(_0197_),
  .ZN(_0198_)
);

NAND3_X1 _1929_ (
  .A1(_0190_),
  .A2(_1119_),
  .A3(_0195_),
  .ZN(_0199_)
);

NAND3_X1 _1930_ (
  .A1(_0198_),
  .A2(_0199_),
  .A3(_0604_),
  .ZN(_0200_)
);

OAI21_X1 _1931_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[15] ),
  .ZN(_0201_)
);

INV_X1 _1932_ (
  .A(_0201_),
  .ZN(_0202_)
);

NAND2_X1 _1933_ (
  .A1(_0200_),
  .A2(_0202_),
  .ZN(_0203_)
);

NAND2_X1 _1934_ (
  .A1(_0387_),
  .A2(result[15]),
  .ZN(_0204_)
);

NAND2_X1 _1935_ (
  .A1(_0203_),
  .A2(_0204_),
  .ZN(_0034_)
);

OAI21_X1 _1936_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[16] ),
  .ZN(_0205_)
);

INV_X1 _1937_ (
  .A(_0205_),
  .ZN(_0206_)
);

NAND2_X1 _1938_ (
  .A1(_1117_),
  .A2(_1119_),
  .ZN(_0207_)
);

NOR2_X1 _1939_ (
  .A1(_0171_),
  .A2(_0207_),
  .ZN(_0208_)
);

NAND3_X1 _1940_ (
  .A1(_0070_),
  .A2(_0130_),
  .A3(_0208_),
  .ZN(_0209_)
);

BUF_X2 _1941_ (
  .A(_1121_),
  .Z(_0210_)
);

INV_X1 _1942_ (
  .A(_1118_),
  .ZN(_0211_)
);

OAI21_X1 _1943_ (
  .A(_0211_),
  .B1(_0197_),
  .B2(_0191_),
  .ZN(_0212_)
);

INV_X1 _1944_ (
  .A(_0212_),
  .ZN(_0213_)
);

OAI21_X1 _1945_ (
  .A(_0213_),
  .B1(_0176_),
  .B2(_0207_),
  .ZN(_0214_)
);

AOI21_X1 _1946_ (
  .A(_0214_),
  .B1(_0208_),
  .B2(_0135_),
  .ZN(_0215_)
);

NAND3_X1 _1947_ (
  .A1(_0209_),
  .A2(_0210_),
  .A3(_0215_),
  .ZN(_0216_)
);

NAND2_X1 _1948_ (
  .A1(_0216_),
  .A2(_0604_),
  .ZN(_0217_)
);

AOI21_X1 _1949_ (
  .A(_0210_),
  .B1(_0209_),
  .B2(_0215_),
  .ZN(_0218_)
);

OAI21_X1 _1950_ (
  .A(_0206_),
  .B1(_0217_),
  .B2(_0218_),
  .ZN(_0219_)
);

NAND2_X1 _1951_ (
  .A1(_0387_),
  .A2(result[16]),
  .ZN(_0220_)
);

NAND2_X1 _1952_ (
  .A1(_0219_),
  .A2(_0220_),
  .ZN(_0035_)
);

OAI21_X1 _1953_ (
  .A(_0371_),
  .B1(_0594_),
  .B2(\ext_mult_res[17] ),
  .ZN(_0221_)
);

INV_X1 _1954_ (
  .A(_0221_),
  .ZN(_0222_)
);

OAI21_X1 _1955_ (
  .A(_0599_),
  .B1(_0589_),
  .B2(_0598_),
  .ZN(_0223_)
);

INV_X1 _1956_ (
  .A(_0223_),
  .ZN(_0224_)
);

OAI21_X1 _1957_ (
  .A(_0622_),
  .B1(_0224_),
  .B2(_0617_),
  .ZN(_0225_)
);

NAND2_X1 _1958_ (
  .A1(_0225_),
  .A2(_0164_),
  .ZN(_0226_)
);

INV_X1 _1959_ (
  .A(_0150_),
  .ZN(_0227_)
);

NAND2_X1 _1960_ (
  .A1(_0226_),
  .A2(_0227_),
  .ZN(_0228_)
);

NAND2_X2 _1961_ (
  .A1(_1119_),
  .A2(_0210_),
  .ZN(_0229_)
);

NOR2_X2 _1962_ (
  .A1(_0188_),
  .A2(_0229_),
  .ZN(_0230_)
);

AND2_X1 _1963_ (
  .A1(_0152_),
  .A2(_0230_),
  .ZN(_0231_)
);

NAND2_X1 _1964_ (
  .A1(_0228_),
  .A2(_0231_),
  .ZN(_0232_)
);

INV_X1 _1965_ (
  .A(_0229_),
  .ZN(_0233_)
);

NAND2_X1 _1966_ (
  .A1(_0192_),
  .A2(_0233_),
  .ZN(_0234_)
);

INV_X1 _1967_ (
  .A(_1120_),
  .ZN(_0235_)
);

INV_X1 _1968_ (
  .A(_0210_),
  .ZN(_0236_)
);

OAI21_X1 _1969_ (
  .A(_0235_),
  .B1(_0236_),
  .B2(_0211_),
  .ZN(_0237_)
);

INV_X1 _1970_ (
  .A(_0237_),
  .ZN(_0238_)
);

NAND2_X1 _1971_ (
  .A1(_0234_),
  .A2(_0238_),
  .ZN(_0239_)
);

AOI21_X1 _1972_ (
  .A(_0239_),
  .B1(_0230_),
  .B2(_0159_),
  .ZN(_0240_)
);

AND3_X1 _1973_ (
  .A1(_0618_),
  .A2(_1091_),
  .A3(_1093_),
  .ZN(_0241_)
);

NAND4_X1 _1974_ (
  .A1(_0231_),
  .A2(_0241_),
  .A3(_0164_),
  .A4(_1088_),
  .ZN(_0242_)
);

NAND3_X1 _1975_ (
  .A1(_0232_),
  .A2(_0240_),
  .A3(_0242_),
  .ZN(_0243_)
);

INV_X1 _1976_ (
  .A(_1123_),
  .ZN(_0244_)
);

NAND2_X1 _1977_ (
  .A1(_0243_),
  .A2(_0244_),
  .ZN(_0245_)
);

NAND2_X1 _1978_ (
  .A1(_0245_),
  .A2(_0604_),
  .ZN(_0246_)
);

NOR2_X1 _1979_ (
  .A1(_0243_),
  .A2(_0244_),
  .ZN(_0247_)
);

OAI21_X1 _1980_ (
  .A(_0222_),
  .B1(_0246_),
  .B2(_0247_),
  .ZN(_0248_)
);

NAND2_X1 _1981_ (
  .A1(_0387_),
  .A2(result[17]),
  .ZN(_0249_)
);

NAND2_X1 _1982_ (
  .A1(_0248_),
  .A2(_0249_),
  .ZN(_0036_)
);

NOR2_X1 _1983_ (
  .A1(_0368_),
  .A2(result[18]),
  .ZN(_0250_)
);

NAND2_X1 _1984_ (
  .A1(_0092_),
  .A2(_0097_),
  .ZN(_0251_)
);

NAND2_X1 _1985_ (
  .A1(_0210_),
  .A2(_1123_),
  .ZN(_0252_)
);

NOR2_X1 _1986_ (
  .A1(_0207_),
  .A2(_0252_),
  .ZN(_0253_)
);

AND2_X1 _1987_ (
  .A1(_0172_),
  .A2(_0253_),
  .ZN(_0254_)
);

NAND2_X1 _1988_ (
  .A1(_0251_),
  .A2(_0254_),
  .ZN(_0255_)
);

INV_X1 _1989_ (
  .A(_1122_),
  .ZN(_0256_)
);

OAI21_X1 _1990_ (
  .A(_0256_),
  .B1(_0244_),
  .B2(_0235_),
  .ZN(_0257_)
);

INV_X1 _1991_ (
  .A(_0257_),
  .ZN(_0258_)
);

OAI21_X1 _1992_ (
  .A(_0258_),
  .B1(_0213_),
  .B2(_0252_),
  .ZN(_0259_)
);

AOI21_X1 _1993_ (
  .A(_0259_),
  .B1(_0253_),
  .B2(_0177_),
  .ZN(_0260_)
);

NAND4_X1 _1994_ (
  .A1(_0254_),
  .A2(_0091_),
  .A3(_0098_),
  .A4(_0099_),
  .ZN(_0261_)
);

NAND3_X1 _1995_ (
  .A1(_0255_),
  .A2(_0260_),
  .A3(_0261_),
  .ZN(_0262_)
);

NAND2_X1 _1996_ (
  .A1(_0262_),
  .A2(_1125_),
  .ZN(_0263_)
);

INV_X1 _1997_ (
  .A(_1125_),
  .ZN(_0264_)
);

NAND4_X1 _1998_ (
  .A1(_0255_),
  .A2(_0260_),
  .A3(_0264_),
  .A4(_0261_),
  .ZN(_0265_)
);

NAND3_X1 _1999_ (
  .A1(_0263_),
  .A2(_0265_),
  .A3(_0584_),
  .ZN(_0266_)
);

NAND2_X1 _2000_ (
  .A1(_0581_),
  .A2(\ext_mult_res[18] ),
  .ZN(_0267_)
);

NAND2_X1 _2001_ (
  .A1(_0267_),
  .A2(_0371_),
  .ZN(_0268_)
);

INV_X1 _2002_ (
  .A(_0268_),
  .ZN(_0269_)
);

AOI21_X1 _2003_ (
  .A(_0250_),
  .B1(_0266_),
  .B2(_0269_),
  .ZN(_0037_)
);

NOR2_X1 _2004_ (
  .A1(_0368_),
  .A2(result[19]),
  .ZN(_0270_)
);

NAND2_X1 _2005_ (
  .A1(_1123_),
  .A2(_1125_),
  .ZN(_0271_)
);

NOR2_X1 _2006_ (
  .A1(_0229_),
  .A2(_0271_),
  .ZN(_0272_)
);

AND2_X1 _2007_ (
  .A1(_0189_),
  .A2(_0272_),
  .ZN(_0273_)
);

NAND2_X1 _2008_ (
  .A1(_0115_),
  .A2(_0273_),
  .ZN(_0274_)
);

INV_X1 _2009_ (
  .A(_1124_),
  .ZN(_0275_)
);

OAI21_X1 _2010_ (
  .A(_0275_),
  .B1(_0264_),
  .B2(_0256_),
  .ZN(_0276_)
);

INV_X1 _2011_ (
  .A(_0276_),
  .ZN(_0277_)
);

OAI21_X1 _2012_ (
  .A(_0277_),
  .B1(_0238_),
  .B2(_0271_),
  .ZN(_0278_)
);

AOI21_X1 _2013_ (
  .A(_0278_),
  .B1(_0272_),
  .B2(_0194_),
  .ZN(_0279_)
);

NAND3_X1 _2014_ (
  .A1(_0118_),
  .A2(_0119_),
  .A3(_0273_),
  .ZN(_0280_)
);

NAND3_X1 _2015_ (
  .A1(_0274_),
  .A2(_0279_),
  .A3(_0280_),
  .ZN(_0281_)
);

NAND2_X1 _2016_ (
  .A1(_0281_),
  .A2(_1127_),
  .ZN(_0282_)
);

INV_X1 _2017_ (
  .A(_1127_),
  .ZN(_0283_)
);

NAND4_X1 _2018_ (
  .A1(_0274_),
  .A2(_0279_),
  .A3(_0283_),
  .A4(_0280_),
  .ZN(_0284_)
);

NAND3_X1 _2019_ (
  .A1(_0282_),
  .A2(_0284_),
  .A3(_0584_),
  .ZN(_0285_)
);

AOI21_X1 _2020_ (
  .A(_0270_),
  .B1(_0285_),
  .B2(_0269_),
  .ZN(_0038_)
);

NOR2_X1 _2021_ (
  .A1(_0368_),
  .A2(result[20]),
  .ZN(_0286_)
);

NAND2_X1 _2022_ (
  .A1(_1125_),
  .A2(_1127_),
  .ZN(_0287_)
);

NOR2_X1 _2023_ (
  .A1(_0252_),
  .A2(_0287_),
  .ZN(_0288_)
);

AND2_X1 _2024_ (
  .A1(_0208_),
  .A2(_0288_),
  .ZN(_0289_)
);

NAND2_X1 _2025_ (
  .A1(_0137_),
  .A2(_0289_),
  .ZN(_0290_)
);

INV_X1 _2026_ (
  .A(_1126_),
  .ZN(_0291_)
);

OAI21_X1 _2027_ (
  .A(_0291_),
  .B1(_0283_),
  .B2(_0275_),
  .ZN(_0292_)
);

INV_X1 _2028_ (
  .A(_0292_),
  .ZN(_0293_)
);

OAI21_X1 _2029_ (
  .A(_0293_),
  .B1(_0258_),
  .B2(_0287_),
  .ZN(_0294_)
);

AOI21_X1 _2030_ (
  .A(_0294_),
  .B1(_0288_),
  .B2(_0214_),
  .ZN(_0295_)
);

NAND3_X1 _2031_ (
  .A1(_0612_),
  .A2(_0140_),
  .A3(_0289_),
  .ZN(_0296_)
);

NAND3_X1 _2032_ (
  .A1(_0290_),
  .A2(_0295_),
  .A3(_0296_),
  .ZN(_0297_)
);

NAND2_X1 _2033_ (
  .A1(_0297_),
  .A2(_1129_),
  .ZN(_0298_)
);

INV_X1 _2034_ (
  .A(_1129_),
  .ZN(_0299_)
);

NAND4_X1 _2035_ (
  .A1(_0290_),
  .A2(_0295_),
  .A3(_0299_),
  .A4(_0296_),
  .ZN(_0300_)
);

NAND3_X1 _2036_ (
  .A1(_0298_),
  .A2(_0300_),
  .A3(_0584_),
  .ZN(_0301_)
);

AOI21_X1 _2037_ (
  .A(_0286_),
  .B1(_0301_),
  .B2(_0269_),
  .ZN(_0039_)
);

NAND2_X1 _2038_ (
  .A1(_1127_),
  .A2(_1129_),
  .ZN(_0302_)
);

NOR2_X1 _2039_ (
  .A1(_0271_),
  .A2(_0302_),
  .ZN(_0303_)
);

NAND2_X1 _2040_ (
  .A1(_0230_),
  .A2(_0303_),
  .ZN(_0304_)
);

INV_X1 _2041_ (
  .A(_0304_),
  .ZN(_0305_)
);

NAND2_X1 _2042_ (
  .A1(_0161_),
  .A2(_0305_),
  .ZN(_0306_)
);

INV_X1 _2043_ (
  .A(_0303_),
  .ZN(_0307_)
);

AOI21_X1 _2044_ (
  .A(_0307_),
  .B1(_0234_),
  .B2(_0238_),
  .ZN(_0308_)
);

INV_X1 _2045_ (
  .A(_1128_),
  .ZN(_0309_)
);

OAI21_X1 _2046_ (
  .A(_0309_),
  .B1(_0299_),
  .B2(_0291_),
  .ZN(_0310_)
);

INV_X1 _2047_ (
  .A(_0310_),
  .ZN(_0311_)
);

OAI21_X1 _2048_ (
  .A(_0311_),
  .B1(_0277_),
  .B2(_0302_),
  .ZN(_0312_)
);

NOR2_X1 _2049_ (
  .A1(_0308_),
  .A2(_0312_),
  .ZN(_0313_)
);

NOR2_X1 _2050_ (
  .A1(_0165_),
  .A2(_0304_),
  .ZN(_0314_)
);

NAND2_X1 _2051_ (
  .A1(_0623_),
  .A2(_0314_),
  .ZN(_0315_)
);

XOR2_X1 _2052_ (
  .A(\ext_mult_res[18] ),
  .B(result[21]),
  .Z(_0316_)
);

NAND4_X1 _2053_ (
  .A1(_0306_),
  .A2(_0313_),
  .A3(_0315_),
  .A4(_0316_),
  .ZN(_0317_)
);

NAND3_X1 _2054_ (
  .A1(_0306_),
  .A2(_0313_),
  .A3(_0315_),
  .ZN(_0318_)
);

INV_X1 _2055_ (
  .A(_0316_),
  .ZN(_0319_)
);

NAND2_X1 _2056_ (
  .A1(_0318_),
  .A2(_0319_),
  .ZN(_0320_)
);

NAND2_X1 _2057_ (
  .A1(_0317_),
  .A2(_0320_),
  .ZN(_0321_)
);

NAND2_X1 _2058_ (
  .A1(_0321_),
  .A2(_0594_),
  .ZN(_0322_)
);

NAND2_X1 _2059_ (
  .A1(_0322_),
  .A2(_0267_),
  .ZN(_0323_)
);

NAND2_X1 _2060_ (
  .A1(_0323_),
  .A2(_0372_),
  .ZN(_0324_)
);

NAND2_X1 _2061_ (
  .A1(_0387_),
  .A2(result[21]),
  .ZN(_0325_)
);

NAND2_X1 _2062_ (
  .A1(_0324_),
  .A2(_0325_),
  .ZN(_0040_)
);

FA_X1 _2063_ (
  .A(_0676_),
  .B(_0677_),
  .CI(_0678_),
  .CO(_0679_),
  .S(_0680_)
);

FA_X1 _2064_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0684_),
  .S(_0685_)
);

FA_X1 _2065_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0689_),
  .S(_0690_)
);

FA_X1 _2066_ (
  .A(_0690_),
  .B(_0684_),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0692_),
  .S(_0693_)
);

FA_X1 _2067_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0697_),
  .S(_0698_)
);

FA_X1 _2068_ (
  .A(_0698_),
  .B(_0699_),
  .CI(_0700_),
  .CO(_0701_),
  .S(_0702_)
);

FA_X1 _2069_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0706_),
  .S(_0707_)
);

FA_X1 _2070_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0711_),
  .S(_0712_)
);

FA_X1 _2071_ (
  .A(_0707_),
  .B(_0697_),
  .CI(_0712_),
  .CO(_0713_),
  .S(_0714_)
);

FA_X1 _2072_ (
  .A(_0715_),
  .B(_0716_),
  .CI(_0717_),
  .CO(_0718_),
  .S(_0719_)
);

FA_X1 _2073_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0723_),
  .S(_0724_)
);

FA_X1 _2074_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0728_),
  .S(_0729_)
);

FA_X1 _2075_ (
  .A(_0724_),
  .B(_0706_),
  .CI(_0729_),
  .CO(_0730_),
  .S(_0731_)
);

FA_X1 _2076_ (
  .A(_0731_),
  .B(_0713_),
  .CI(_0732_),
  .CO(_0733_),
  .S(_0734_)
);

FA_X1 _2077_ (
  .A(_0735_),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0738_),
  .S(_0739_)
);

FA_X1 _2078_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0743_),
  .S(_0744_)
);

FA_X1 _2079_ (
  .A(_0744_),
  .B(_0739_),
  .CI(_0745_),
  .CO(_0746_),
  .S(_0747_)
);

FA_X1 _2080_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0751_),
  .S(_0752_)
);

FA_X1 _2081_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0756_),
  .S(_0757_)
);

FA_X1 _2082_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0761_),
  .S(_0762_)
);

FA_X1 _2083_ (
  .A(_0765_),
  .B(_0766_),
  .CI(_0767_),
  .CO(_0768_),
  .S(_0769_)
);

FA_X1 _2084_ (
  .A(_0770_),
  .B(_0747_),
  .CI(_0771_),
  .CO(_0772_),
  .S(_0773_)
);

FA_X1 _2085_ (
  .A(_0757_),
  .B(_0774_),
  .CI(_0775_),
  .CO(_0776_),
  .S(_0777_)
);

FA_X1 _2086_ (
  .A(_0778_),
  .B(_0779_),
  .CI(_0780_),
  .CO(_0781_),
  .S(_0782_)
);

FA_X1 _2087_ (
  .A(_0777_),
  .B(_0730_),
  .CI(_0784_),
  .CO(_0783_),
  .S(_0785_)
);

FA_X1 _2088_ (
  .A(_0786_),
  .B(_0733_),
  .CI(_0787_),
  .CO(_0788_),
  .S(_0789_)
);

FA_X1 _2089_ (
  .A(_0790_),
  .B(_0791_),
  .CI(_0792_),
  .CO(_0793_),
  .S(_0794_)
);

FA_X1 _2090_ (
  .A(_0795_),
  .B(_0796_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0798_),
  .S(_0799_)
);

FA_X1 _2091_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0803_),
  .S(_0804_)
);

FA_X1 _2092_ (
  .A(_0799_),
  .B(_0738_),
  .CI(_0804_),
  .CO(_0805_),
  .S(_0806_)
);

FA_X1 _2093_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0809_),
  .S(_0810_)
);

FA_X1 _2094_ (
  .A(_0811_),
  .B(_0812_),
  .CI(_0813_),
  .CO(_0814_),
  .S(_0815_)
);

FA_X1 _2095_ (
  .A(_0806_),
  .B(_0746_),
  .CI(_0815_),
  .CO(_0816_),
  .S(_0817_)
);

FA_X1 _2096_ (
  .A(_0817_),
  .B(_0772_),
  .CI(_0818_),
  .CO(_0819_),
  .S(_0820_)
);

FA_X1 _2097_ (
  .A(_0821_),
  .B(_0822_),
  .CI(_0823_),
  .CO(_0824_),
  .S(_0825_)
);

FA_X1 _2098_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0829_),
  .S(_0830_)
);

FA_X1 _2099_ (
  .A(_0825_),
  .B(_0798_),
  .CI(_0830_),
  .CO(_0831_),
  .S(_0832_)
);

FA_X1 _2100_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0835_),
  .S(_0836_)
);

FA_X1 _2101_ (
  .A(_0837_),
  .B(_0838_),
  .CI(_0839_),
  .CO(_0840_),
  .S(_0841_)
);

FA_X1 _2102_ (
  .A(_0841_),
  .B(_0832_),
  .CI(_0805_),
  .CO(_0842_),
  .S(_0843_)
);

FA_X1 _2103_ (
  .A(_0816_),
  .B(_0843_),
  .CI(_0844_),
  .CO(_0845_),
  .S(_0846_)
);

FA_X1 _2104_ (
  .A(_0847_),
  .B(_0848_),
  .CI(_0849_),
  .CO(_0850_),
  .S(_0851_)
);

FA_X1 _2105_ (
  .A(_0852_),
  .B(_0853_),
  .CI(_0854_),
  .CO(_0855_),
  .S(_0856_)
);

FA_X1 _2106_ (
  .A(_0857_),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0860_),
  .S(_0861_)
);

FA_X1 _2107_ (
  .A(_0862_),
  .B(_0824_),
  .CI(_0861_),
  .CO(_0863_),
  .S(_0864_)
);

FA_X1 _2108_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0867_),
  .S(_0868_)
);

FA_X1 _2109_ (
  .A(_0829_),
  .B(_0868_),
  .CI(_0835_),
  .CO(_0869_),
  .S(_0870_)
);

FA_X1 _2110_ (
  .A(_0864_),
  .B(_0831_),
  .CI(_0870_),
  .CO(_0871_),
  .S(_0872_)
);

FA_X1 _2111_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0874_),
  .S(_0875_)
);

FA_X1 _2112_ (
  .A(_0872_),
  .B(_0842_),
  .CI(_0876_),
  .CO(_0877_),
  .S(_0878_)
);

FA_X1 _2113_ (
  .A(_0878_),
  .B(_0845_),
  .CI(_0879_),
  .CO(_0880_),
  .S(_0881_)
);

FA_X1 _2114_ (
  .A(_0852_),
  .B(_0882_),
  .CI(_0854_),
  .CO(_0883_),
  .S(_0884_)
);

FA_X1 _2115_ (
  .A(_0885_),
  .B(_0886_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0888_),
  .S(_0889_)
);

FA_X1 _2116_ (
  .A(_0890_),
  .B(_0891_),
  .CI(_0889_),
  .CO(_0892_),
  .S(_0893_)
);

FA_X1 _2117_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0896_),
  .S(_0897_)
);

FA_X1 _2118_ (
  .A(_0860_),
  .B(_0897_),
  .CI(_0867_),
  .CO(_0898_),
  .S(_0899_)
);

FA_X1 _2119_ (
  .A(_0893_),
  .B(_0863_),
  .CI(_0899_),
  .CO(_0900_),
  .S(_0901_)
);

FA_X1 _2120_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0902_),
  .S(_0903_)
);

FA_X1 _2121_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(_0904_),
  .CI(_0905_),
  .CO(_0906_),
  .S(_0907_)
);

FA_X1 _2122_ (
  .A(_0908_),
  .B(_0909_),
  .CI(_0910_),
  .CO(_0911_),
  .S(_0912_)
);

FA_X1 _2123_ (
  .A(_0901_),
  .B(_0871_),
  .CI(_0913_),
  .CO(_0914_),
  .S(_0915_)
);

FA_X1 _2124_ (
  .A(_0915_),
  .B(_0877_),
  .CI(_0916_),
  .CO(_0917_),
  .S(_0918_)
);

FA_X1 _2125_ (
  .A(_0919_),
  .B(_0920_),
  .CI(_0921_),
  .CO(_0922_),
  .S(_0923_)
);

FA_X1 _2126_ (
  .A(_0924_),
  .B(_0923_),
  .CI(_0890_),
  .CO(_0925_),
  .S(_0926_)
);

FA_X1 _2127_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0929_),
  .S(_0930_)
);

FA_X1 _2128_ (
  .A(_0888_),
  .B(_0930_),
  .CI(_0896_),
  .CO(_0931_),
  .S(_0932_)
);

FA_X1 _2129_ (
  .A(_0926_),
  .B(_0892_),
  .CI(_0932_),
  .CO(_0933_),
  .S(_0934_)
);

FA_X1 _2130_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0935_),
  .S(_0936_)
);

FA_X1 _2131_ (
  .A(_0937_),
  .B(_0938_),
  .CI(_0902_),
  .CO(_0939_),
  .S(_0940_)
);

FA_X1 _2132_ (
  .A(_0898_),
  .B(_0940_),
  .CI(_0906_),
  .CO(_0943_),
  .S(_0944_)
);

FA_X1 _2133_ (
  .A(_0934_),
  .B(_0900_),
  .CI(_0944_),
  .CO(_0945_),
  .S(_0946_)
);

FA_X1 _2134_ (
  .A(_0947_),
  .B(_0948_),
  .CI(_0911_),
  .CO(_0949_),
  .S(_0950_)
);

FA_X1 _2135_ (
  .A(_0951_),
  .B(_0952_),
  .CI(_0953_),
  .CO(_0954_),
  .S(_0955_)
);

FA_X1 _2136_ (
  .A(_0924_),
  .B(_0956_),
  .CI(_0890_),
  .CO(_0957_),
  .S(_0958_)
);

FA_X1 _2137_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(_0959_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0961_),
  .S(_0962_)
);

FA_X1 _2138_ (
  .A(_0922_),
  .B(_0962_),
  .CI(_0929_),
  .CO(_0963_),
  .S(_0964_)
);

FA_X1 _2139_ (
  .A(_0958_),
  .B(_0925_),
  .CI(_0964_),
  .CO(_0965_),
  .S(_0966_)
);

FA_X1 _2140_ (
  .A(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0967_),
  .S(_0968_)
);

FA_X1 _2141_ (
  .A(_0969_),
  .B(_0970_),
  .CI(_0935_),
  .CO(_0971_),
  .S(_0972_)
);

FA_X1 _2142_ (
  .A(_0974_),
  .B(_0975_),
  .CI(_0976_),
  .CO(_0977_),
  .S(_0978_)
);

FA_X1 _2143_ (
  .A(_0966_),
  .B(_0933_),
  .CI(_0978_),
  .CO(_0979_),
  .S(_0980_)
);

FA_X1 _2144_ (
  .A(_0981_),
  .B(_0982_),
  .CI(_0983_),
  .CO(_0984_),
  .S(_0985_)
);

FA_X1 _2145_ (
  .A(_0951_),
  .B(_0986_),
  .CI(_0952_),
  .CO(_0987_),
  .S(_0988_)
);

FA_X1 _2146_ (
  .A(_0924_),
  .B(_0989_),
  .CI(_0890_),
  .CO(_0990_),
  .S(_0991_)
);

FA_X1 _2147_ (
  .A(_0992_),
  .B(_0993_),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0994_),
  .S(_0995_)
);

FA_X1 _2148_ (
  .A(_0995_),
  .B(_0961_),
  .CI(_0996_),
  .CO(_0997_),
  .S(_0998_)
);

FA_X1 _2149_ (
  .A(_0998_),
  .B(_0991_),
  .CI(_0957_),
  .CO(_0999_),
  .S(_1000_)
);

FA_X1 _2150_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_1004_),
  .S(_1005_)
);

FA_X1 _2151_ (
  .A(_1005_),
  .B(_1006_),
  .CI(_0903_),
  .CO(_1007_),
  .S(_1008_)
);

FA_X1 _2152_ (
  .A(_1009_),
  .B(_1008_),
  .CI(_1010_),
  .CO(_1011_),
  .S(_1012_)
);

FA_X1 _2153_ (
  .A(_1000_),
  .B(_0965_),
  .CI(_1012_),
  .CO(_1013_),
  .S(_1014_)
);

FA_X1 _2154_ (
  .A(_1014_),
  .B(_0979_),
  .CI(_1015_),
  .CO(_1016_),
  .S(_1017_)
);

FA_X1 _2155_ (
  .A(_1018_),
  .B(_0984_),
  .CI(_1019_),
  .CO(_1020_),
  .S(_1021_)
);

FA_X1 _2156_ (
  .A(_1022_),
  .B(_1023_),
  .CI(_1024_),
  .CO(_1025_),
  .S(_1026_)
);

FA_X1 _2157_ (
  .A(_1027_),
  .B(_1028_),
  .CI(_0994_),
  .CO(_1029_),
  .S(_1030_)
);

FA_X1 _2158_ (
  .A(_0990_),
  .B(_1030_),
  .CI(_0991_),
  .CO(_1031_),
  .S(_1032_)
);

FA_X1 _2159_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_1034_),
  .S(_1035_)
);

FA_X1 _2160_ (
  .A(_1035_),
  .B(_1004_),
  .CI(_0936_),
  .CO(_1036_),
  .S(_1037_)
);

FA_X1 _2161_ (
  .A(_0997_),
  .B(_1038_),
  .CI(_1039_),
  .CO(_1040_),
  .S(_1041_)
);

FA_X1 _2162_ (
  .A(_1032_),
  .B(_0999_),
  .CI(_1041_),
  .CO(_1042_),
  .S(_1043_)
);

FA_X1 _2163_ (
  .A(_1043_),
  .B(_1013_),
  .CI(_1044_),
  .CO(_1045_),
  .S(_1046_)
);

FA_X1 _2164_ (
  .A(_1047_),
  .B(_1048_),
  .CI(_1049_),
  .CO(_1050_),
  .S(_1051_)
);

FA_X1 _2165_ (
  .A(_1052_),
  .B(_1053_),
  .CI(_1054_),
  .CO(_1055_),
  .S(_1056_)
);

FA_X1 _2166_ (
  .A(_1027_),
  .B(_1057_),
  .CI(_1058_),
  .CO(_1059_),
  .S(_1060_)
);

FA_X1 _2167_ (
  .A(_0990_),
  .B(_1060_),
  .CI(_0991_),
  .CO(_1061_),
  .S(_1062_)
);

FA_X1 _2168_ (
  .A(_0993_),
  .B(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CI(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_1063_),
  .S(_1064_)
);

FA_X1 _2169_ (
  .A(_1034_),
  .B(_1064_),
  .CI(_0968_),
  .CO(_1065_),
  .S(_1066_)
);

FA_X1 _2170_ (
  .A(_1066_),
  .B(_1036_),
  .CI(_1067_),
  .CO(_1068_),
  .S(_1069_)
);

FA_X1 _2171_ (
  .A(_1069_),
  .B(_1062_),
  .CI(_1031_),
  .CO(_1070_),
  .S(_1071_)
);

FA_X1 _2172_ (
  .A(_0973_),
  .B(_0875_),
  .CI(_1072_),
  .CO(_1073_),
  .S(_1074_)
);

FA_X1 _2173_ (
  .A(_1075_),
  .B(_1076_),
  .CI(_1077_),
  .CO(_1078_),
  .S(_1079_)
);

FA_X1 _2174_ (
  .A(_1071_),
  .B(_1042_),
  .CI(_1080_),
  .CO(_1081_),
  .S(_1082_)
);

FA_X1 _2175_ (
  .A(_1083_),
  .B(_1084_),
  .CI(_1085_),
  .CO(_1086_),
  .S(_1087_)
);

HA_X1 _2176_ (
  .A(result[0]),
  .B(\ext_mult_res[0] ),
  .CO(_1088_),
  .S(_1089_)
);

HA_X1 _2177_ (
  .A(result[1]),
  .B(\ext_mult_res[1] ),
  .CO(_1090_),
  .S(_1091_)
);

HA_X1 _2178_ (
  .A(result[2]),
  .B(\ext_mult_res[2] ),
  .CO(_1092_),
  .S(_1093_)
);

HA_X1 _2179_ (
  .A(result[3]),
  .B(\ext_mult_res[3] ),
  .CO(_1094_),
  .S(_1095_)
);

HA_X1 _2180_ (
  .A(result[4]),
  .B(\ext_mult_res[4] ),
  .CO(_1096_),
  .S(_1097_)
);

HA_X1 _2181_ (
  .A(result[5]),
  .B(\ext_mult_res[5] ),
  .CO(_1098_),
  .S(_1099_)
);

HA_X1 _2182_ (
  .A(result[6]),
  .B(\ext_mult_res[6] ),
  .CO(_1100_),
  .S(_1101_)
);

HA_X1 _2183_ (
  .A(result[7]),
  .B(\ext_mult_res[7] ),
  .CO(_1102_),
  .S(_1103_)
);

HA_X1 _2184_ (
  .A(result[8]),
  .B(\ext_mult_res[8] ),
  .CO(_1104_),
  .S(_1105_)
);

HA_X1 _2185_ (
  .A(result[9]),
  .B(\ext_mult_res[9] ),
  .CO(_1106_),
  .S(_1107_)
);

HA_X1 _2186_ (
  .A(result[10]),
  .B(\ext_mult_res[10] ),
  .CO(_1108_),
  .S(_1109_)
);

HA_X1 _2187_ (
  .A(result[11]),
  .B(\ext_mult_res[11] ),
  .CO(_1110_),
  .S(_1111_)
);

HA_X1 _2188_ (
  .A(result[12]),
  .B(\ext_mult_res[12] ),
  .CO(_1112_),
  .S(_1113_)
);

HA_X1 _2189_ (
  .A(result[13]),
  .B(\ext_mult_res[13] ),
  .CO(_1114_),
  .S(_1115_)
);

HA_X1 _2190_ (
  .A(result[14]),
  .B(\ext_mult_res[14] ),
  .CO(_1116_),
  .S(_1117_)
);

HA_X1 _2191_ (
  .A(result[15]),
  .B(\ext_mult_res[15] ),
  .CO(_1118_),
  .S(_1119_)
);

HA_X1 _2192_ (
  .A(result[16]),
  .B(\ext_mult_res[16] ),
  .CO(_1120_),
  .S(_1121_)
);

HA_X1 _2193_ (
  .A(result[17]),
  .B(\ext_mult_res[17] ),
  .CO(_1122_),
  .S(_1123_)
);

HA_X1 _2194_ (
  .A(result[18]),
  .B(\ext_mult_res[18] ),
  .CO(_1124_),
  .S(_1125_)
);

HA_X1 _2195_ (
  .A(result[19]),
  .B(\ext_mult_res[18] ),
  .CO(_1126_),
  .S(_1127_)
);

HA_X1 _2196_ (
  .A(result[20]),
  .B(\ext_mult_res[18] ),
  .CO(_1128_),
  .S(_1129_)
);

HA_X1 _2197_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_1132_),
  .S(_1133_)
);

HA_X1 _2198_ (
  .A(_0685_),
  .B(_1132_),
  .CO(_1134_),
  .S(_1135_)
);

HA_X1 _2199_ (
  .A(_0693_),
  .B(_1134_),
  .CO(_1136_),
  .S(_1137_)
);

HA_X1 _2200_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0717_),
  .S(_1140_)
);

HA_X1 _2201_ (
  .A(_1141_),
  .B(_0692_),
  .CO(_1142_),
  .S(_1143_)
);

HA_X1 _2202_ (
  .A(_1143_),
  .B(_1136_),
  .CO(_1144_),
  .S(_1145_)
);

HA_X1 _2203_ (
  .A(_0719_),
  .B(_1142_),
  .CO(_1146_),
  .S(_1147_)
);

HA_X1 _2204_ (
  .A(_1147_),
  .B(_1144_),
  .CO(_1148_),
  .S(_1149_)
);

HA_X1 _2205_ (
  .A(_1150_),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_1152_),
  .S(_1153_)
);

HA_X1 _2206_ (
  .A(_1154_),
  .B(_0718_),
  .CO(_1155_),
  .S(_1156_)
);

HA_X1 _2207_ (
  .A(_1156_),
  .B(_1146_),
  .CO(_1157_),
  .S(_1158_)
);

HA_X1 _2208_ (
  .A(_1158_),
  .B(_1148_),
  .CO(_1159_),
  .S(_1160_)
);

HA_X1 _2209_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_0767_),
  .S(_1162_)
);

HA_X1 _2210_ (
  .A(_1163_),
  .B(_1162_),
  .CO(_0780_),
  .S(_1164_)
);

HA_X1 _2211_ (
  .A(_0782_),
  .B(_1165_),
  .CO(_1166_),
  .S(_1167_)
);

HA_X1 _2212_ (
  .A(_1167_),
  .B(_1168_),
  .CO(_1169_),
  .S(_1170_)
);

HA_X1 _2213_ (
  .A(_1171_),
  .B(_1155_),
  .CO(_1168_),
  .S(_1172_)
);

HA_X1 _2214_ (
  .A(_1170_),
  .B(_1173_),
  .CO(_1174_),
  .S(_1175_)
);

HA_X1 _2215_ (
  .A(_1172_),
  .B(_1157_),
  .CO(_1173_),
  .S(_1176_)
);

HA_X1 _2216_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(_0768_),
  .CO(_0847_),
  .S(_1178_)
);

HA_X1 _2217_ (
  .A(_1179_),
  .B(_0781_),
  .CO(_1180_),
  .S(_1181_)
);

HA_X1 _2218_ (
  .A(_1181_),
  .B(_1166_),
  .CO(_1182_),
  .S(_1183_)
);

HA_X1 _2219_ (
  .A(_1183_),
  .B(_1169_),
  .CO(_1184_),
  .S(_1185_)
);

HA_X1 _2220_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .CO(_1072_),
  .S(_0941_)
);

HA_X1 _2221_ (
  .A(_0814_),
  .B(_0941_),
  .CO(_1186_),
  .S(_1187_)
);

HA_X1 _2222_ (
  .A(_0851_),
  .B(_1180_),
  .CO(_1188_),
  .S(_1189_)
);

HA_X1 _2223_ (
  .A(_1189_),
  .B(_1182_),
  .CO(_1190_),
  .S(_1191_)
);

HA_X1 _2224_ (
  .A(_0875_),
  .B(_1072_),
  .CO(_0910_),
  .S(_1192_)
);

HA_X1 _2225_ (
  .A(_0840_),
  .B(_1192_),
  .CO(_1193_),
  .S(_1194_)
);

HA_X1 _2226_ (
  .A(_0881_),
  .B(_0850_),
  .CO(_1195_),
  .S(_1196_)
);

HA_X1 _2227_ (
  .A(_1196_),
  .B(_1188_),
  .CO(_1197_),
  .S(_1198_)
);

HA_X1 _2228_ (
  .A(_1199_),
  .B(_0918_),
  .CO(_1200_),
  .S(_1201_)
);

HA_X1 _2229_ (
  .A(_1195_),
  .B(_1201_),
  .CO(_1202_),
  .S(_1203_)
);

HA_X1 _2230_ (
  .A(_1204_),
  .B(_1205_),
  .CO(_1206_),
  .S(_1207_)
);

HA_X1 _2231_ (
  .A(_1207_),
  .B(_1200_),
  .CO(_1208_),
  .S(_1209_)
);

HA_X1 _2232_ (
  .A(_1210_),
  .B(_1072_),
  .CO(_1019_),
  .S(_0981_)
);

HA_X1 _2233_ (
  .A(_1211_),
  .B(_0949_),
  .CO(_1212_),
  .S(_1213_)
);

HA_X1 _2234_ (
  .A(_1213_),
  .B(_1206_),
  .CO(_1214_),
  .S(_1215_)
);

HA_X1 _2235_ (
  .A(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 ),
  .B(_0874_),
  .CO(_1217_),
  .S(_1218_)
);

HA_X1 _2236_ (
  .A(_0977_),
  .B(_1218_),
  .CO(_1049_),
  .S(_1219_)
);

HA_X1 _2237_ (
  .A(_1021_),
  .B(_1212_),
  .CO(_1220_),
  .S(_1221_)
);

HA_X1 _2238_ (
  .A(_1222_),
  .B(_1216_),
  .CO(_1223_),
  .S(_1224_)
);

HA_X1 _2239_ (
  .A(_0941_),
  .B(_0942_),
  .CO(_1225_),
  .S(_1226_)
);

HA_X1 _2240_ (
  .A(_1226_),
  .B(_1217_),
  .CO(_1077_),
  .S(_1227_)
);

HA_X1 _2241_ (
  .A(_1011_),
  .B(_1227_),
  .CO(_1085_),
  .S(_1228_)
);

HA_X1 _2242_ (
  .A(_1051_),
  .B(_1020_),
  .CO(_1229_),
  .S(_1230_)
);

HA_X1 _2243_ (
  .A(_1074_),
  .B(_1225_),
  .CO(_1231_),
  .S(_1076_)
);

HA_X1 _2244_ (
  .A(_1087_),
  .B(_1050_),
  .CO(_1232_),
  .S(_1233_)
);

HA_X1 _2245_ (
  .A(_1176_),
  .B(_1159_),
  .CO(_1177_),
  .S(_1234_)
);

DFF_X1 \ext_mult_res[0]$_DFFE_PP_  (
  .D(_0000_),
  .CK(clk),
  .Q(\ext_mult_res[0] ),
  .QN(_0675_)
);

DFF_X1 \ext_mult_res[10]$_DFFE_PP_  (
  .D(_0010_),
  .CK(clk),
  .Q(\ext_mult_res[10] ),
  .QN(_0666_)
);

DFF_X1 \ext_mult_res[11]$_DFFE_PP_  (
  .D(_0011_),
  .CK(clk),
  .Q(\ext_mult_res[11] ),
  .QN(_0665_)
);

DFF_X1 \ext_mult_res[12]$_DFFE_PP_  (
  .D(_0012_),
  .CK(clk),
  .Q(\ext_mult_res[12] ),
  .QN(_0664_)
);

DFF_X1 \ext_mult_res[13]$_DFFE_PP_  (
  .D(_0013_),
  .CK(clk),
  .Q(\ext_mult_res[13] ),
  .QN(_0663_)
);

DFF_X1 \ext_mult_res[14]$_DFFE_PP_  (
  .D(_0014_),
  .CK(clk),
  .Q(\ext_mult_res[14] ),
  .QN(_0662_)
);

DFF_X1 \ext_mult_res[15]$_DFFE_PP_  (
  .D(_0015_),
  .CK(clk),
  .Q(\ext_mult_res[15] ),
  .QN(_0661_)
);

DFF_X1 \ext_mult_res[16]$_DFFE_PP_  (
  .D(_0016_),
  .CK(clk),
  .Q(\ext_mult_res[16] ),
  .QN(_0660_)
);

DFF_X1 \ext_mult_res[17]$_DFFE_PP_  (
  .D(_0017_),
  .CK(clk),
  .Q(\ext_mult_res[17] ),
  .QN(_0659_)
);

DFF_X1 \ext_mult_res[1]$_DFFE_PP_  (
  .D(_0001_),
  .CK(clk),
  .Q(\ext_mult_res[1] ),
  .QN(_0677_)
);

DFF_X1 \ext_mult_res[21]$_DFFE_PP_  (
  .D(_0018_),
  .CK(clk),
  .Q(\ext_mult_res[18] ),
  .QN(_0658_)
);

DFF_X1 \ext_mult_res[2]$_DFFE_PP_  (
  .D(_0002_),
  .CK(clk),
  .Q(\ext_mult_res[2] ),
  .QN(_0674_)
);

DFF_X1 \ext_mult_res[3]$_DFFE_PP_  (
  .D(_0003_),
  .CK(clk),
  .Q(\ext_mult_res[3] ),
  .QN(_0673_)
);

DFF_X1 \ext_mult_res[4]$_DFFE_PP_  (
  .D(_0004_),
  .CK(clk),
  .Q(\ext_mult_res[4] ),
  .QN(_0672_)
);

DFF_X1 \ext_mult_res[5]$_DFFE_PP_  (
  .D(_0005_),
  .CK(clk),
  .Q(\ext_mult_res[5] ),
  .QN(_0671_)
);

DFF_X1 \ext_mult_res[6]$_DFFE_PP_  (
  .D(_0006_),
  .CK(clk),
  .Q(\ext_mult_res[6] ),
  .QN(_0670_)
);

DFF_X1 \ext_mult_res[7]$_DFFE_PP_  (
  .D(_0007_),
  .CK(clk),
  .Q(\ext_mult_res[7] ),
  .QN(_0669_)
);

DFF_X1 \ext_mult_res[8]$_DFFE_PP_  (
  .D(_0008_),
  .CK(clk),
  .Q(\ext_mult_res[8] ),
  .QN(_0668_)
);

DFF_X1 \ext_mult_res[9]$_DFFE_PP_  (
  .D(_0009_),
  .CK(clk),
  .Q(\ext_mult_res[9] ),
  .QN(_0667_)
);

DFF_X1 \result[0]$_DFFE_PP_  (
  .D(_0019_),
  .CK(clk),
  .Q(result[0]),
  .QN(_0657_)
);

DFF_X1 \result[10]$_DFFE_PP_  (
  .D(_0029_),
  .CK(clk),
  .Q(result[10]),
  .QN(_0648_)
);

DFF_X1 \result[11]$_DFFE_PP_  (
  .D(_0030_),
  .CK(clk),
  .Q(result[11]),
  .QN(_0647_)
);

DFF_X1 \result[12]$_DFFE_PP_  (
  .D(_0031_),
  .CK(clk),
  .Q(result[12]),
  .QN(_0646_)
);

DFF_X1 \result[13]$_DFFE_PP_  (
  .D(_0032_),
  .CK(clk),
  .Q(result[13]),
  .QN(_0645_)
);

DFF_X1 \result[14]$_DFFE_PP_  (
  .D(_0033_),
  .CK(clk),
  .Q(result[14]),
  .QN(_0644_)
);

DFF_X1 \result[15]$_DFFE_PP_  (
  .D(_0034_),
  .CK(clk),
  .Q(result[15]),
  .QN(_0643_)
);

DFF_X1 \result[16]$_DFFE_PP_  (
  .D(_0035_),
  .CK(clk),
  .Q(result[16]),
  .QN(_0642_)
);

DFF_X1 \result[17]$_DFFE_PP_  (
  .D(_0036_),
  .CK(clk),
  .Q(result[17]),
  .QN(_0641_)
);

DFF_X1 \result[18]$_DFFE_PP_  (
  .D(_0037_),
  .CK(clk),
  .Q(result[18]),
  .QN(_0640_)
);

DFF_X1 \result[19]$_DFFE_PP_  (
  .D(_0038_),
  .CK(clk),
  .Q(result[19]),
  .QN(_0639_)
);

DFF_X1 \result[1]$_DFFE_PP_  (
  .D(_0020_),
  .CK(clk),
  .Q(result[1]),
  .QN(_0676_)
);

DFF_X1 \result[20]$_DFFE_PP_  (
  .D(_0039_),
  .CK(clk),
  .Q(result[20]),
  .QN(_0638_)
);

DFF_X1 \result[21]$_DFFE_PP_  (
  .D(_0040_),
  .CK(clk),
  .Q(result[21]),
  .QN(_0637_)
);

DFF_X1 \result[2]$_DFFE_PP_  (
  .D(_0021_),
  .CK(clk),
  .Q(result[2]),
  .QN(_0656_)
);

DFF_X1 \result[3]$_DFFE_PP_  (
  .D(_0022_),
  .CK(clk),
  .Q(result[3]),
  .QN(_0655_)
);

DFF_X1 \result[4]$_DFFE_PP_  (
  .D(_0023_),
  .CK(clk),
  .Q(result[4]),
  .QN(_0654_)
);

DFF_X1 \result[5]$_DFFE_PP_  (
  .D(_0024_),
  .CK(clk),
  .Q(result[5]),
  .QN(_0653_)
);

DFF_X1 \result[6]$_DFFE_PP_  (
  .D(_0025_),
  .CK(clk),
  .Q(result[6]),
  .QN(_0652_)
);

DFF_X1 \result[7]$_DFFE_PP_  (
  .D(_0026_),
  .CK(clk),
  .Q(result[7]),
  .QN(_0651_)
);

DFF_X1 \result[8]$_DFFE_PP_  (
  .D(_0027_),
  .CK(clk),
  .Q(result[8]),
  .QN(_0650_)
);

DFF_X1 \result[9]$_DFFE_PP_  (
  .D(_0028_),
  .CK(clk),
  .Q(result[9]),
  .QN(_0649_)
);

LOGIC0_X1 \logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644  (
  .Z(\logic0_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 )
);

LOGIC1_X1 \logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644  (
  .Z(\logic1_naja_$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644 )
);

INV_X1 _1283__reduced (
  .A(_0326_),
  .ZN(_0735_)
);

INV_X1 _1308__reduced (
  .A(_0333_),
  .ZN(_0796_)
);

INV_X1 _1319__reduced (
  .A(_0339_),
  .ZN(_0823_)
);

INV_X1 _1328__reduced (
  .A(_0341_),
  .ZN(_0857_)
);

INV_X1 _1337__reduced (
  .A(_0354_),
  .ZN(_0886_)
);

INV_X1 _1345__reduced (
  .A(_0355_),
  .ZN(_0921_)
);

INV_X1 _1353__reduced (
  .A(_0348_),
  .ZN(_0959_)
);

INV_X1 _1359__reduced (
  .A(din[7]),
  .ZN(_0993_)
);

NOR2_X1 _1473__reduced (
  .A1(_0370_),
  .A2(_0372_),
  .ZN(_0000_)
);

INV_X1 _1634__reduced (
  .A(_0993_),
  .ZN(_0516_)
);

INV_X1 _1636__reduced (
  .A(_0516_),
  .ZN(_0518_)
);

NAND2_X1 _1638__reduced (
  .A1(_0516_),
  .A2(_0358_),
  .ZN(_0520_)
);

NAND2_X1 _1643__reduced (
  .A1(_0516_),
  .A2(_0524_),
  .ZN(_0525_)
);

NAND2_X1 _1662__reduced (
  .A1(_0540_),
  .A2(_0541_),
  .ZN(_0544_)
);

INV_X1 _1663__reduced (
  .A(_0544_),
  .ZN(_0545_)
);

NAND2_X1 _1667__reduced (
  .A1(_0544_),
  .A2(_0546_),
  .ZN(_0549_)
);
endmodule //$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644

module \$paramod$04fdc4f446e06e0744e44efd615d1158fec3aeb8\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _197_ (
  .A(x[1]),
  .ZN(_180_)
);

INV_X1 _198_ (
  .A(x[0]),
  .ZN(_179_)
);

BUF_X1 _199_ (
  .A(ena),
  .Z(_110_)
);

BUF_X2 _200_ (
  .A(_110_),
  .Z(_111_)
);

NOR2_X1 _201_ (
  .A1(\coef[10] ),
  .A2(_111_),
  .ZN(_112_)
);

BUF_X4 _202_ (
  .A(x[2]),
  .Z(_113_)
);

INV_X8 _203_ (
  .A(_113_),
  .ZN(_114_)
);

NAND2_X1 _204_ (
  .A1(_114_),
  .A2(_181_),
  .ZN(_115_)
);

INV_X1 _205_ (
  .A(_195_),
  .ZN(_116_)
);

BUF_X8 _206_ (
  .A(_113_),
  .Z(_117_)
);

NAND2_X2 _207_ (
  .A1(_116_),
  .A2(_117_),
  .ZN(_118_)
);

BUF_X8 _208_ (
  .A(y[0]),
  .Z(_119_)
);

INV_X8 _209_ (
  .A(_119_),
  .ZN(_120_)
);

BUF_X16 _210_ (
  .A(_120_),
  .Z(_121_)
);

NAND3_X1 _211_ (
  .A1(_115_),
  .A2(_118_),
  .A3(_121_),
  .ZN(_122_)
);

NAND2_X1 _212_ (
  .A1(_114_),
  .A2(_116_),
  .ZN(_123_)
);

NAND2_X2 _213_ (
  .A1(_117_),
  .A2(_181_),
  .ZN(_124_)
);

NAND3_X1 _214_ (
  .A1(_123_),
  .A2(_119_),
  .A3(_124_),
  .ZN(_125_)
);

NAND2_X1 _215_ (
  .A1(_122_),
  .A2(_125_),
  .ZN(_126_)
);

BUF_X4 _216_ (
  .A(y[2]),
  .Z(_127_)
);

INV_X4 _217_ (
  .A(_127_),
  .ZN(_128_)
);

BUF_X4 _218_ (
  .A(y[1]),
  .Z(_129_)
);

NAND2_X1 _219_ (
  .A1(_128_),
  .A2(_129_),
  .ZN(_130_)
);

INV_X1 _220_ (
  .A(_130_),
  .ZN(_131_)
);

NAND2_X1 _221_ (
  .A1(_126_),
  .A2(_131_),
  .ZN(_132_)
);

NAND2_X1 _222_ (
  .A1(_114_),
  .A2(_193_),
  .ZN(_133_)
);

INV_X1 _223_ (
  .A(_183_),
  .ZN(_134_)
);

NAND2_X2 _224_ (
  .A1(_134_),
  .A2(_117_),
  .ZN(_135_)
);

NAND3_X1 _225_ (
  .A1(_133_),
  .A2(_135_),
  .A3(_121_),
  .ZN(_136_)
);

NAND2_X1 _226_ (
  .A1(_114_),
  .A2(_134_),
  .ZN(_137_)
);

BUF_X4 _227_ (
  .A(_119_),
  .Z(_138_)
);

NAND2_X2 _228_ (
  .A1(_117_),
  .A2(_193_),
  .ZN(_139_)
);

NAND3_X1 _229_ (
  .A1(_137_),
  .A2(_138_),
  .A3(_139_),
  .ZN(_140_)
);

NAND2_X1 _230_ (
  .A1(_136_),
  .A2(_140_),
  .ZN(_141_)
);

NOR2_X4 _231_ (
  .A1(_128_),
  .A2(_129_),
  .ZN(_142_)
);

NAND2_X1 _232_ (
  .A1(_141_),
  .A2(_142_),
  .ZN(_143_)
);

NAND2_X1 _233_ (
  .A1(_132_),
  .A2(_143_),
  .ZN(_144_)
);

NAND2_X1 _234_ (
  .A1(_129_),
  .A2(_127_),
  .ZN(_145_)
);

OR2_X2 _235_ (
  .A1(_191_),
  .A2(_117_),
  .ZN(_146_)
);

NAND2_X1 _236_ (
  .A1(_117_),
  .A2(_185_),
  .ZN(_147_)
);

NAND3_X1 _237_ (
  .A1(_146_),
  .A2(_138_),
  .A3(_147_),
  .ZN(_148_)
);

OR2_X2 _238_ (
  .A1(_187_),
  .A2(_113_),
  .ZN(_149_)
);

NAND2_X2 _239_ (
  .A1(_117_),
  .A2(_189_),
  .ZN(_150_)
);

NAND3_X1 _240_ (
  .A1(_149_),
  .A2(_121_),
  .A3(_150_),
  .ZN(_151_)
);

AOI21_X1 _241_ (
  .A(_145_),
  .B1(_148_),
  .B2(_151_),
  .ZN(_152_)
);

NOR2_X2 _242_ (
  .A1(_144_),
  .A2(_152_),
  .ZN(_153_)
);

INV_X1 _243_ (
  .A(_110_),
  .ZN(_154_)
);

INV_X1 _244_ (
  .A(_189_),
  .ZN(_155_)
);

NAND2_X1 _245_ (
  .A1(_114_),
  .A2(_155_),
  .ZN(_156_)
);

NAND2_X1 _246_ (
  .A1(_117_),
  .A2(_187_),
  .ZN(_157_)
);

NAND2_X1 _247_ (
  .A1(_156_),
  .A2(_157_),
  .ZN(_158_)
);

NAND2_X1 _248_ (
  .A1(_158_),
  .A2(_121_),
  .ZN(_159_)
);

INV_X1 _249_ (
  .A(_185_),
  .ZN(_160_)
);

NAND2_X1 _250_ (
  .A1(_114_),
  .A2(_160_),
  .ZN(_161_)
);

NAND2_X1 _251_ (
  .A1(_113_),
  .A2(_191_),
  .ZN(_162_)
);

NAND2_X1 _252_ (
  .A1(_161_),
  .A2(_162_),
  .ZN(_163_)
);

NAND2_X1 _253_ (
  .A1(_163_),
  .A2(_138_),
  .ZN(_164_)
);

NAND2_X1 _254_ (
  .A1(_159_),
  .A2(_164_),
  .ZN(_165_)
);

INV_X4 _255_ (
  .A(_129_),
  .ZN(_166_)
);

NAND2_X2 _256_ (
  .A1(_166_),
  .A2(_128_),
  .ZN(_167_)
);

INV_X2 _257_ (
  .A(_167_),
  .ZN(_168_)
);

AOI21_X1 _258_ (
  .A(_154_),
  .B1(_165_),
  .B2(_168_),
  .ZN(_169_)
);

AOI21_X2 _259_ (
  .A(_112_),
  .B1(_153_),
  .B2(_169_),
  .ZN(_000_)
);

NAND2_X4 _260_ (
  .A1(_117_),
  .A2(_119_),
  .ZN(_009_)
);

NAND2_X1 _261_ (
  .A1(_009_),
  .A2(_166_),
  .ZN(_010_)
);

INV_X1 _262_ (
  .A(_010_),
  .ZN(_011_)
);

NAND2_X1 _263_ (
  .A1(_151_),
  .A2(_011_),
  .ZN(_012_)
);

NAND3_X1 _264_ (
  .A1(_133_),
  .A2(_135_),
  .A3(_138_),
  .ZN(_013_)
);

OAI21_X1 _265_ (
  .A(_129_),
  .B1(_179_),
  .B2(_119_),
  .ZN(_014_)
);

INV_X1 _266_ (
  .A(_014_),
  .ZN(_015_)
);

NAND2_X1 _267_ (
  .A1(_013_),
  .A2(_015_),
  .ZN(_016_)
);

NAND3_X1 _268_ (
  .A1(_012_),
  .A2(_016_),
  .A3(_127_),
  .ZN(_017_)
);

AOI21_X4 _269_ (
  .A(_166_),
  .B1(_120_),
  .B2(_114_),
  .ZN(_018_)
);

NAND2_X1 _270_ (
  .A1(_164_),
  .A2(_018_),
  .ZN(_019_)
);

NAND3_X1 _271_ (
  .A1(_123_),
  .A2(_121_),
  .A3(_124_),
  .ZN(_020_)
);

AOI21_X1 _272_ (
  .A(_129_),
  .B1(_179_),
  .B2(_138_),
  .ZN(_021_)
);

NAND2_X1 _273_ (
  .A1(_020_),
  .A2(_021_),
  .ZN(_022_)
);

NAND3_X1 _274_ (
  .A1(_019_),
  .A2(_022_),
  .A3(_128_),
  .ZN(_023_)
);

NAND2_X1 _275_ (
  .A1(_017_),
  .A2(_023_),
  .ZN(_024_)
);

NAND2_X1 _276_ (
  .A1(_024_),
  .A2(_111_),
  .ZN(_025_)
);

NAND2_X1 _277_ (
  .A1(_154_),
  .A2(\coef[21] ),
  .ZN(_026_)
);

NAND2_X1 _278_ (
  .A1(_025_),
  .A2(_026_),
  .ZN(_001_)
);

NOR2_X1 _279_ (
  .A1(_111_),
  .A2(\coef[23] ),
  .ZN(_027_)
);

NAND2_X1 _280_ (
  .A1(_119_),
  .A2(x[0]),
  .ZN(_028_)
);

OAI21_X1 _281_ (
  .A(_028_),
  .B1(_117_),
  .B2(_119_),
  .ZN(_029_)
);

AND2_X1 _282_ (
  .A1(_029_),
  .A2(_168_),
  .ZN(_030_)
);

NAND2_X2 _283_ (
  .A1(_149_),
  .A2(_150_),
  .ZN(_031_)
);

NOR2_X1 _284_ (
  .A1(_031_),
  .A2(_130_),
  .ZN(_032_)
);

AND2_X1 _285_ (
  .A1(_163_),
  .A2(_142_),
  .ZN(_033_)
);

NOR3_X1 _286_ (
  .A1(_030_),
  .A2(_032_),
  .A3(_033_),
  .ZN(_034_)
);

NAND2_X4 _287_ (
  .A1(_121_),
  .A2(_179_),
  .ZN(_035_)
);

NAND2_X2 _288_ (
  .A1(_035_),
  .A2(_009_),
  .ZN(_036_)
);

INV_X1 _289_ (
  .A(_145_),
  .ZN(_037_)
);

AOI21_X1 _290_ (
  .A(_154_),
  .B1(_036_),
  .B2(_037_),
  .ZN(_038_)
);

AOI21_X1 _291_ (
  .A(_027_),
  .B1(_034_),
  .B2(_038_),
  .ZN(_002_)
);

NOR2_X1 _292_ (
  .A1(_111_),
  .A2(\coef[24] ),
  .ZN(_039_)
);

NAND3_X2 _293_ (
  .A1(_115_),
  .A2(_118_),
  .A3(_119_),
  .ZN(_040_)
);

INV_X1 _294_ (
  .A(_182_),
  .ZN(_041_)
);

NAND2_X2 _295_ (
  .A1(_114_),
  .A2(_041_),
  .ZN(_042_)
);

NAND2_X1 _296_ (
  .A1(_113_),
  .A2(_182_),
  .ZN(_043_)
);

NAND3_X2 _297_ (
  .A1(_042_),
  .A2(_121_),
  .A3(_043_),
  .ZN(_044_)
);

NAND2_X1 _298_ (
  .A1(_040_),
  .A2(_044_),
  .ZN(_045_)
);

NAND2_X1 _299_ (
  .A1(_045_),
  .A2(_168_),
  .ZN(_046_)
);

NAND2_X1 _300_ (
  .A1(_042_),
  .A2(_043_),
  .ZN(_047_)
);

NAND2_X1 _301_ (
  .A1(_047_),
  .A2(_138_),
  .ZN(_048_)
);

NAND3_X2 _302_ (
  .A1(_137_),
  .A2(_121_),
  .A3(_139_),
  .ZN(_049_)
);

NAND2_X1 _303_ (
  .A1(_048_),
  .A2(_049_),
  .ZN(_050_)
);

INV_X1 _304_ (
  .A(_050_),
  .ZN(_051_)
);

OAI21_X1 _305_ (
  .A(_046_),
  .B1(_051_),
  .B2(_145_),
  .ZN(_052_)
);

INV_X1 _306_ (
  .A(_052_),
  .ZN(_053_)
);

NAND3_X1 _307_ (
  .A1(_161_),
  .A2(_121_),
  .A3(_162_),
  .ZN(_054_)
);

NAND3_X1 _308_ (
  .A1(_054_),
  .A2(_127_),
  .A3(_011_),
  .ZN(_055_)
);

NAND2_X1 _309_ (
  .A1(_055_),
  .A2(_111_),
  .ZN(_056_)
);

NAND2_X2 _310_ (
  .A1(_031_),
  .A2(_138_),
  .ZN(_057_)
);

NAND2_X1 _311_ (
  .A1(_057_),
  .A2(_018_),
  .ZN(_058_)
);

NOR2_X1 _312_ (
  .A1(_058_),
  .A2(_127_),
  .ZN(_059_)
);

NOR2_X1 _313_ (
  .A1(_056_),
  .A2(_059_),
  .ZN(_060_)
);

AOI21_X2 _314_ (
  .A(_039_),
  .B1(_053_),
  .B2(_060_),
  .ZN(_003_)
);

NOR2_X1 _315_ (
  .A1(_111_),
  .A2(\coef[26] ),
  .ZN(_061_)
);

NAND2_X1 _316_ (
  .A1(_020_),
  .A2(_028_),
  .ZN(_062_)
);

NAND2_X1 _317_ (
  .A1(_062_),
  .A2(_166_),
  .ZN(_063_)
);

NAND3_X1 _318_ (
  .A1(_054_),
  .A2(_129_),
  .A3(_028_),
  .ZN(_064_)
);

NAND2_X1 _319_ (
  .A1(_063_),
  .A2(_064_),
  .ZN(_065_)
);

NAND2_X1 _320_ (
  .A1(_065_),
  .A2(_127_),
  .ZN(_066_)
);

AND2_X2 _321_ (
  .A1(_168_),
  .A2(_035_),
  .ZN(_067_)
);

NAND2_X1 _322_ (
  .A1(_057_),
  .A2(_067_),
  .ZN(_068_)
);

NAND2_X1 _323_ (
  .A1(_068_),
  .A2(_111_),
  .ZN(_069_)
);

AOI21_X1 _324_ (
  .A(_130_),
  .B1(_013_),
  .B2(_035_),
  .ZN(_070_)
);

NOR2_X2 _325_ (
  .A1(_069_),
  .A2(_070_),
  .ZN(_071_)
);

AOI21_X2 _326_ (
  .A(_061_),
  .B1(_066_),
  .B2(_071_),
  .ZN(_004_)
);

NOR2_X1 _327_ (
  .A1(_111_),
  .A2(\coef[13] ),
  .ZN(_072_)
);

NAND3_X1 _328_ (
  .A1(_156_),
  .A2(_138_),
  .A3(_157_),
  .ZN(_073_)
);

NAND3_X1 _329_ (
  .A1(_044_),
  .A2(_073_),
  .A3(_037_),
  .ZN(_074_)
);

NAND2_X1 _330_ (
  .A1(_119_),
  .A2(x[1]),
  .ZN(_075_)
);

NAND2_X1 _331_ (
  .A1(_049_),
  .A2(_075_),
  .ZN(_076_)
);

NAND2_X1 _332_ (
  .A1(_076_),
  .A2(_142_),
  .ZN(_077_)
);

NAND2_X1 _333_ (
  .A1(_074_),
  .A2(_077_),
  .ZN(_078_)
);

NAND2_X1 _334_ (
  .A1(_048_),
  .A2(_168_),
  .ZN(_079_)
);

AOI21_X1 _335_ (
  .A(_138_),
  .B1(_146_),
  .B2(_147_),
  .ZN(_080_)
);

NOR2_X1 _336_ (
  .A1(_079_),
  .A2(_080_),
  .ZN(_081_)
);

NOR2_X2 _337_ (
  .A1(_078_),
  .A2(_081_),
  .ZN(_082_)
);

NAND2_X4 _338_ (
  .A1(_121_),
  .A2(_180_),
  .ZN(_083_)
);

NAND2_X1 _339_ (
  .A1(_040_),
  .A2(_083_),
  .ZN(_084_)
);

AOI21_X1 _340_ (
  .A(_154_),
  .B1(_084_),
  .B2(_131_),
  .ZN(_085_)
);

AOI21_X2 _341_ (
  .A(_072_),
  .B1(_082_),
  .B2(_085_),
  .ZN(_005_)
);

OR2_X1 _342_ (
  .A1(\coef[28] ),
  .A2(_110_),
  .ZN(_086_)
);

INV_X1 _343_ (
  .A(_142_),
  .ZN(_087_)
);

OAI21_X2 _344_ (
  .A(_110_),
  .B1(_036_),
  .B2(_087_),
  .ZN(_088_)
);

NOR2_X1 _345_ (
  .A1(_029_),
  .A2(_130_),
  .ZN(_089_)
);

NOR2_X2 _346_ (
  .A1(_088_),
  .A2(_089_),
  .ZN(_090_)
);

NAND2_X1 _347_ (
  .A1(_048_),
  .A2(_083_),
  .ZN(_091_)
);

NAND2_X1 _348_ (
  .A1(_091_),
  .A2(_037_),
  .ZN(_092_)
);

NAND2_X1 _349_ (
  .A1(_090_),
  .A2(_092_),
  .ZN(_093_)
);

AOI21_X1 _350_ (
  .A(_167_),
  .B1(_044_),
  .B2(_075_),
  .ZN(_094_)
);

OAI21_X1 _351_ (
  .A(_086_),
  .B1(_093_),
  .B2(_094_),
  .ZN(_095_)
);

INV_X1 _352_ (
  .A(_095_),
  .ZN(_006_)
);

OR2_X1 _353_ (
  .A1(\coef[29] ),
  .A2(_110_),
  .ZN(_096_)
);

NAND2_X1 _354_ (
  .A1(_018_),
  .A2(_075_),
  .ZN(_097_)
);

NOR2_X1 _355_ (
  .A1(_097_),
  .A2(_127_),
  .ZN(_098_)
);

NAND3_X2 _356_ (
  .A1(_142_),
  .A2(_083_),
  .A3(_009_),
  .ZN(_099_)
);

NAND2_X2 _357_ (
  .A1(_099_),
  .A2(_110_),
  .ZN(_100_)
);

NOR2_X2 _358_ (
  .A1(_098_),
  .A2(_100_),
  .ZN(_101_)
);

NAND2_X1 _359_ (
  .A1(_136_),
  .A2(_040_),
  .ZN(_102_)
);

NAND2_X1 _360_ (
  .A1(_102_),
  .A2(_037_),
  .ZN(_103_)
);

NAND2_X1 _361_ (
  .A1(_101_),
  .A2(_103_),
  .ZN(_104_)
);

AOI21_X1 _362_ (
  .A(_167_),
  .B1(_125_),
  .B2(_049_),
  .ZN(_105_)
);

OAI21_X1 _363_ (
  .A(_096_),
  .B1(_104_),
  .B2(_105_),
  .ZN(_106_)
);

INV_X1 _364_ (
  .A(_106_),
  .ZN(_007_)
);

NOR2_X1 _365_ (
  .A1(_111_),
  .A2(\coef[30] ),
  .ZN(_107_)
);

OAI21_X1 _366_ (
  .A(_130_),
  .B1(_142_),
  .B2(_138_),
  .ZN(_108_)
);

XNOR2_X1 _367_ (
  .A(_108_),
  .B(_114_),
  .ZN(_109_)
);

AOI21_X1 _368_ (
  .A(_107_),
  .B1(_109_),
  .B2(_111_),
  .ZN(_008_)
);

HA_X1 _369_ (
  .A(_179_),
  .B(_180_),
  .CO(_181_),
  .S(_182_)
);

HA_X1 _370_ (
  .A(_179_),
  .B(_180_),
  .CO(_183_),
  .S(_184_)
);

HA_X1 _371_ (
  .A(_179_),
  .B(x[1]),
  .CO(_185_),
  .S(_186_)
);

HA_X1 _372_ (
  .A(_179_),
  .B(x[1]),
  .CO(_187_),
  .S(_188_)
);

HA_X1 _373_ (
  .A(x[0]),
  .B(_180_),
  .CO(_189_),
  .S(_190_)
);

HA_X1 _374_ (
  .A(x[0]),
  .B(_180_),
  .CO(_191_),
  .S(_192_)
);

HA_X1 _375_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_193_),
  .S(_194_)
);

HA_X1 _376_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_195_),
  .S(_196_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_177_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_176_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_175_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_178_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_174_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_173_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_172_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_171_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_170_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$04fdc4f446e06e0744e44efd615d1158fec3aeb8\dctu

module \$paramod$fa85f450a22557b2687ca86acb15721a7fddf8e7\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

CLKBUF_X3 _067_ (
  .A(ena),
  .Z(_008_)
);

NOR2_X1 _068_ (
  .A1(\coef[21] ),
  .A2(_008_),
  .ZN(_009_)
);

INV_X1 _069_ (
  .A(_008_),
  .ZN(_010_)
);

INV_X2 _070_ (
  .A(x[0]),
  .ZN(_011_)
);

NAND2_X1 _071_ (
  .A1(_011_),
  .A2(x[1]),
  .ZN(_012_)
);

INV_X2 _072_ (
  .A(x[1]),
  .ZN(_013_)
);

NAND2_X1 _073_ (
  .A1(_013_),
  .A2(x[0]),
  .ZN(_014_)
);

NAND2_X4 _074_ (
  .A1(_012_),
  .A2(_014_),
  .ZN(_015_)
);

NAND2_X2 _075_ (
  .A1(_015_),
  .A2(y[0]),
  .ZN(_016_)
);

NAND2_X2 _076_ (
  .A1(_013_),
  .A2(_011_),
  .ZN(_017_)
);

NAND2_X1 _077_ (
  .A1(x[1]),
  .A2(x[0]),
  .ZN(_018_)
);

NAND2_X2 _078_ (
  .A1(_017_),
  .A2(_018_),
  .ZN(_019_)
);

INV_X1 _079_ (
  .A(y[0]),
  .ZN(_020_)
);

NAND2_X2 _080_ (
  .A1(_019_),
  .A2(_020_),
  .ZN(_021_)
);

CLKBUF_X3 _081_ (
  .A(y[1]),
  .Z(_022_)
);

INV_X1 _082_ (
  .A(_022_),
  .ZN(_023_)
);

NAND3_X2 _083_ (
  .A1(_016_),
  .A2(_021_),
  .A3(_023_),
  .ZN(_024_)
);

NAND2_X4 _084_ (
  .A1(_015_),
  .A2(_022_),
  .ZN(_025_)
);

INV_X2 _085_ (
  .A(_025_),
  .ZN(_026_)
);

BUF_X1 _086_ (
  .A(y[2]),
  .Z(_027_)
);

INV_X1 _087_ (
  .A(_027_),
  .ZN(_028_)
);

NOR2_X1 _088_ (
  .A1(_026_),
  .A2(_028_),
  .ZN(_029_)
);

AOI21_X1 _089_ (
  .A(_010_),
  .B1(_024_),
  .B2(_029_),
  .ZN(_030_)
);

NAND3_X2 _090_ (
  .A1(_016_),
  .A2(_021_),
  .A3(_022_),
  .ZN(_031_)
);

NOR2_X4 _091_ (
  .A1(_015_),
  .A2(_022_),
  .ZN(_032_)
);

NOR2_X1 _092_ (
  .A1(_032_),
  .A2(_027_),
  .ZN(_033_)
);

NAND2_X1 _093_ (
  .A1(_031_),
  .A2(_033_),
  .ZN(_034_)
);

AOI21_X2 _094_ (
  .A(_009_),
  .B1(_030_),
  .B2(_034_),
  .ZN(_000_)
);

NOR3_X2 _095_ (
  .A1(_026_),
  .A2(_032_),
  .A3(_010_),
  .ZN(_035_)
);

INV_X1 _096_ (
  .A(\coef[22] ),
  .ZN(_036_)
);

AOI21_X1 _097_ (
  .A(_035_),
  .B1(_036_),
  .B2(_010_),
  .ZN(_001_)
);

NOR2_X1 _098_ (
  .A1(_008_),
  .A2(\coef[23] ),
  .ZN(_037_)
);

XNOR2_X1 _099_ (
  .A(_019_),
  .B(_027_),
  .ZN(_038_)
);

AOI21_X1 _100_ (
  .A(_037_),
  .B1(_038_),
  .B2(_008_),
  .ZN(_002_)
);

INV_X1 _101_ (
  .A(_035_),
  .ZN(_039_)
);

INV_X1 _102_ (
  .A(\coef[14] ),
  .ZN(_040_)
);

OAI21_X1 _103_ (
  .A(_039_),
  .B1(_008_),
  .B2(_040_),
  .ZN(_003_)
);

NAND2_X2 _104_ (
  .A1(_019_),
  .A2(y[0]),
  .ZN(_041_)
);

NAND3_X1 _105_ (
  .A1(_017_),
  .A2(_020_),
  .A3(_018_),
  .ZN(_042_)
);

NAND3_X2 _106_ (
  .A1(_041_),
  .A2(_042_),
  .A3(_022_),
  .ZN(_043_)
);

NOR2_X1 _107_ (
  .A1(_032_),
  .A2(_028_),
  .ZN(_044_)
);

AOI21_X2 _108_ (
  .A(_010_),
  .B1(_043_),
  .B2(_044_),
  .ZN(_045_)
);

NAND3_X2 _109_ (
  .A1(_041_),
  .A2(_042_),
  .A3(_023_),
  .ZN(_046_)
);

NAND3_X1 _110_ (
  .A1(_046_),
  .A2(_028_),
  .A3(_025_),
  .ZN(_047_)
);

NAND2_X1 _111_ (
  .A1(_045_),
  .A2(_047_),
  .ZN(_048_)
);

NAND2_X1 _112_ (
  .A1(_010_),
  .A2(\coef[13] ),
  .ZN(_049_)
);

NAND2_X1 _113_ (
  .A1(_048_),
  .A2(_049_),
  .ZN(_004_)
);

NOR2_X1 _114_ (
  .A1(_008_),
  .A2(\coef[28] ),
  .ZN(_050_)
);

AOI21_X1 _115_ (
  .A(_010_),
  .B1(_043_),
  .B2(_033_),
  .ZN(_051_)
);

NAND3_X1 _116_ (
  .A1(_046_),
  .A2(_027_),
  .A3(_025_),
  .ZN(_052_)
);

AOI21_X2 _117_ (
  .A(_050_),
  .B1(_051_),
  .B2(_052_),
  .ZN(_005_)
);

NAND3_X1 _118_ (
  .A1(_024_),
  .A2(_043_),
  .A3(_028_),
  .ZN(_053_)
);

NAND3_X1 _119_ (
  .A1(_031_),
  .A2(_046_),
  .A3(_027_),
  .ZN(_054_)
);

NAND3_X1 _120_ (
  .A1(_053_),
  .A2(_054_),
  .A3(_008_),
  .ZN(_055_)
);

NAND2_X1 _121_ (
  .A1(_010_),
  .A2(\coef[15] ),
  .ZN(_056_)
);

NAND2_X1 _122_ (
  .A1(_055_),
  .A2(_056_),
  .ZN(_006_)
);

NAND3_X1 _123_ (
  .A1(_016_),
  .A2(_021_),
  .A3(_008_),
  .ZN(_057_)
);

INV_X1 _124_ (
  .A(\coef[12] ),
  .ZN(_058_)
);

OAI21_X1 _125_ (
  .A(_057_),
  .B1(_008_),
  .B2(_058_),
  .ZN(_007_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_066_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_065_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_064_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_063_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_062_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_061_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_060_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_059_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$fa85f450a22557b2687ca86acb15721a7fddf8e7\dctu

module \$paramod$26ce9ce45d1136272d6a188b0b22329681d6199b\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

BUF_X4 _122_ (
  .A(x[2]),
  .Z(_044_)
);

INV_X4 _123_ (
  .A(_044_),
  .ZN(_045_)
);

NAND2_X2 _124_ (
  .A1(_045_),
  .A2(x[0]),
  .ZN(_046_)
);

INV_X1 _125_ (
  .A(x[0]),
  .ZN(_047_)
);

NAND2_X1 _126_ (
  .A1(_047_),
  .A2(_044_),
  .ZN(_048_)
);

NAND2_X2 _127_ (
  .A1(_046_),
  .A2(_048_),
  .ZN(_049_)
);

BUF_X4 _128_ (
  .A(y[0]),
  .Z(_050_)
);

NAND2_X4 _129_ (
  .A1(_049_),
  .A2(_050_),
  .ZN(_051_)
);

INV_X2 _130_ (
  .A(x[1]),
  .ZN(_052_)
);

NAND2_X2 _131_ (
  .A1(_052_),
  .A2(_044_),
  .ZN(_053_)
);

NAND2_X4 _132_ (
  .A1(_045_),
  .A2(x[1]),
  .ZN(_054_)
);

INV_X2 _133_ (
  .A(_050_),
  .ZN(_055_)
);

NAND3_X2 _134_ (
  .A1(_053_),
  .A2(_054_),
  .A3(_055_),
  .ZN(_056_)
);

BUF_X4 _135_ (
  .A(y[1]),
  .Z(_057_)
);

INV_X4 _136_ (
  .A(_057_),
  .ZN(_058_)
);

NAND3_X2 _137_ (
  .A1(_051_),
  .A2(_056_),
  .A3(_058_),
  .ZN(_059_)
);

NAND2_X2 _138_ (
  .A1(_045_),
  .A2(_052_),
  .ZN(_060_)
);

NAND2_X1 _139_ (
  .A1(_044_),
  .A2(x[1]),
  .ZN(_061_)
);

NAND3_X2 _140_ (
  .A1(_060_),
  .A2(_055_),
  .A3(_061_),
  .ZN(_062_)
);

NAND3_X1 _141_ (
  .A1(_051_),
  .A2(_062_),
  .A3(_057_),
  .ZN(_063_)
);

NAND2_X1 _142_ (
  .A1(_059_),
  .A2(_063_),
  .ZN(_064_)
);

BUF_X2 _143_ (
  .A(y[2]),
  .Z(_065_)
);

INV_X1 _144_ (
  .A(_065_),
  .ZN(_066_)
);

NAND2_X1 _145_ (
  .A1(_064_),
  .A2(_066_),
  .ZN(_067_)
);

NAND2_X2 _146_ (
  .A1(_045_),
  .A2(_047_),
  .ZN(_068_)
);

NAND2_X2 _147_ (
  .A1(_044_),
  .A2(x[0]),
  .ZN(_069_)
);

NAND3_X4 _148_ (
  .A1(_068_),
  .A2(_055_),
  .A3(_069_),
  .ZN(_070_)
);

NAND3_X1 _149_ (
  .A1(_060_),
  .A2(_050_),
  .A3(_061_),
  .ZN(_071_)
);

BUF_X4 _150_ (
  .A(_058_),
  .Z(_072_)
);

NAND3_X1 _151_ (
  .A1(_070_),
  .A2(_071_),
  .A3(_072_),
  .ZN(_073_)
);

NAND3_X4 _152_ (
  .A1(_053_),
  .A2(_054_),
  .A3(_050_),
  .ZN(_074_)
);

NAND3_X2 _153_ (
  .A1(_074_),
  .A2(_070_),
  .A3(_057_),
  .ZN(_075_)
);

NAND3_X1 _154_ (
  .A1(_073_),
  .A2(_075_),
  .A3(_065_),
  .ZN(_076_)
);

NAND2_X1 _155_ (
  .A1(_067_),
  .A2(_076_),
  .ZN(_077_)
);

BUF_X1 _156_ (
  .A(ena),
  .Z(_078_)
);

BUF_X2 _157_ (
  .A(_078_),
  .Z(_079_)
);

NAND2_X1 _158_ (
  .A1(_077_),
  .A2(_079_),
  .ZN(_080_)
);

INV_X1 _159_ (
  .A(_078_),
  .ZN(_081_)
);

NAND2_X1 _160_ (
  .A1(_081_),
  .A2(\coef[21] ),
  .ZN(_082_)
);

NAND2_X1 _161_ (
  .A1(_080_),
  .A2(_082_),
  .ZN(_000_)
);

NAND3_X4 _162_ (
  .A1(_074_),
  .A2(_062_),
  .A3(_058_),
  .ZN(_083_)
);

NAND2_X2 _163_ (
  .A1(_053_),
  .A2(_054_),
  .ZN(_084_)
);

NOR2_X2 _164_ (
  .A1(_084_),
  .A2(_072_),
  .ZN(_085_)
);

NOR2_X1 _165_ (
  .A1(_085_),
  .A2(_065_),
  .ZN(_086_)
);

AOI21_X1 _166_ (
  .A(_081_),
  .B1(_083_),
  .B2(_086_),
  .ZN(_087_)
);

NAND3_X1 _167_ (
  .A1(_074_),
  .A2(_062_),
  .A3(_057_),
  .ZN(_088_)
);

NAND2_X1 _168_ (
  .A1(_084_),
  .A2(_072_),
  .ZN(_089_)
);

NAND3_X1 _169_ (
  .A1(_088_),
  .A2(_065_),
  .A3(_089_),
  .ZN(_090_)
);

NAND2_X1 _170_ (
  .A1(_087_),
  .A2(_090_),
  .ZN(_091_)
);

INV_X1 _171_ (
  .A(\coef[22] ),
  .ZN(_092_)
);

OAI21_X1 _172_ (
  .A(_091_),
  .B1(_079_),
  .B2(_092_),
  .ZN(_001_)
);

NOR2_X1 _173_ (
  .A1(_079_),
  .A2(\coef[23] ),
  .ZN(_093_)
);

NAND2_X1 _174_ (
  .A1(_074_),
  .A2(_070_),
  .ZN(_094_)
);

NAND2_X1 _175_ (
  .A1(_094_),
  .A2(_072_),
  .ZN(_095_)
);

AOI21_X1 _176_ (
  .A(_066_),
  .B1(_049_),
  .B2(_057_),
  .ZN(_096_)
);

AOI21_X1 _177_ (
  .A(_081_),
  .B1(_095_),
  .B2(_096_),
  .ZN(_097_)
);

NAND3_X1 _178_ (
  .A1(_051_),
  .A2(_056_),
  .A3(_057_),
  .ZN(_098_)
);

NAND2_X2 _179_ (
  .A1(_068_),
  .A2(_069_),
  .ZN(_099_)
);

AOI21_X1 _180_ (
  .A(_065_),
  .B1(_099_),
  .B2(_072_),
  .ZN(_100_)
);

NAND2_X1 _181_ (
  .A1(_098_),
  .A2(_100_),
  .ZN(_101_)
);

AOI21_X1 _182_ (
  .A(_093_),
  .B1(_097_),
  .B2(_101_),
  .ZN(_002_)
);

NAND3_X2 _183_ (
  .A1(_056_),
  .A2(_071_),
  .A3(_057_),
  .ZN(_102_)
);

NAND2_X1 _184_ (
  .A1(_102_),
  .A2(_083_),
  .ZN(_103_)
);

NAND2_X1 _185_ (
  .A1(_103_),
  .A2(_066_),
  .ZN(_104_)
);

NAND3_X1 _186_ (
  .A1(_102_),
  .A2(_083_),
  .A3(_065_),
  .ZN(_105_)
);

NAND3_X1 _187_ (
  .A1(_104_),
  .A2(_105_),
  .A3(_079_),
  .ZN(_106_)
);

NAND2_X1 _188_ (
  .A1(_081_),
  .A2(\coef[24] ),
  .ZN(_107_)
);

NAND2_X1 _189_ (
  .A1(_106_),
  .A2(_107_),
  .ZN(_003_)
);

NAND2_X1 _190_ (
  .A1(_049_),
  .A2(_072_),
  .ZN(_108_)
);

NAND3_X1 _191_ (
  .A1(_098_),
  .A2(_065_),
  .A3(_108_),
  .ZN(_109_)
);

NOR2_X1 _192_ (
  .A1(_049_),
  .A2(_072_),
  .ZN(_110_)
);

INV_X1 _193_ (
  .A(_110_),
  .ZN(_111_)
);

NAND3_X1 _194_ (
  .A1(_095_),
  .A2(_066_),
  .A3(_111_),
  .ZN(_010_)
);

NAND3_X1 _195_ (
  .A1(_109_),
  .A2(_010_),
  .A3(_079_),
  .ZN(_011_)
);

NAND2_X1 _196_ (
  .A1(_081_),
  .A2(\coef[25] ),
  .ZN(_012_)
);

NAND2_X1 _197_ (
  .A1(_011_),
  .A2(_012_),
  .ZN(_004_)
);

NAND2_X1 _198_ (
  .A1(_075_),
  .A2(_083_),
  .ZN(_013_)
);

NAND2_X1 _199_ (
  .A1(_013_),
  .A2(_066_),
  .ZN(_014_)
);

NAND3_X1 _200_ (
  .A1(_059_),
  .A2(_102_),
  .A3(_065_),
  .ZN(_015_)
);

NAND2_X1 _201_ (
  .A1(_014_),
  .A2(_015_),
  .ZN(_016_)
);

NAND2_X1 _202_ (
  .A1(_016_),
  .A2(_079_),
  .ZN(_017_)
);

NAND2_X1 _203_ (
  .A1(_081_),
  .A2(\coef[26] ),
  .ZN(_018_)
);

NAND2_X1 _204_ (
  .A1(_017_),
  .A2(_018_),
  .ZN(_005_)
);

NAND2_X1 _205_ (
  .A1(_070_),
  .A2(_071_),
  .ZN(_019_)
);

NAND2_X1 _206_ (
  .A1(_019_),
  .A2(_057_),
  .ZN(_020_)
);

NAND3_X1 _207_ (
  .A1(_020_),
  .A2(_095_),
  .A3(_066_),
  .ZN(_021_)
);

NAND3_X1 _208_ (
  .A1(_051_),
  .A2(_062_),
  .A3(_072_),
  .ZN(_022_)
);

NAND3_X1 _209_ (
  .A1(_098_),
  .A2(_022_),
  .A3(_065_),
  .ZN(_023_)
);

NAND3_X1 _210_ (
  .A1(_021_),
  .A2(_023_),
  .A3(_079_),
  .ZN(_024_)
);

NAND2_X1 _211_ (
  .A1(_081_),
  .A2(\coef[27] ),
  .ZN(_025_)
);

NAND2_X1 _212_ (
  .A1(_024_),
  .A2(_025_),
  .ZN(_006_)
);

NAND2_X1 _213_ (
  .A1(_099_),
  .A2(_050_),
  .ZN(_026_)
);

NAND2_X2 _214_ (
  .A1(_026_),
  .A2(_070_),
  .ZN(_027_)
);

NAND2_X1 _215_ (
  .A1(_027_),
  .A2(_057_),
  .ZN(_028_)
);

NAND2_X1 _216_ (
  .A1(_028_),
  .A2(_100_),
  .ZN(_029_)
);

NAND2_X1 _217_ (
  .A1(_027_),
  .A2(_072_),
  .ZN(_030_)
);

NAND2_X1 _218_ (
  .A1(_030_),
  .A2(_096_),
  .ZN(_031_)
);

NAND3_X1 _219_ (
  .A1(_029_),
  .A2(_031_),
  .A3(_079_),
  .ZN(_032_)
);

INV_X1 _220_ (
  .A(\coef[28] ),
  .ZN(_033_)
);

OAI21_X1 _221_ (
  .A(_032_),
  .B1(_079_),
  .B2(_033_),
  .ZN(_007_)
);

NOR2_X1 _222_ (
  .A1(_078_),
  .A2(\coef[15] ),
  .ZN(_034_)
);

INV_X1 _223_ (
  .A(_059_),
  .ZN(_035_)
);

OAI21_X1 _224_ (
  .A(_066_),
  .B1(_035_),
  .B2(_085_),
  .ZN(_036_)
);

INV_X1 _225_ (
  .A(_084_),
  .ZN(_037_)
);

AOI21_X1 _226_ (
  .A(_066_),
  .B1(_037_),
  .B2(_072_),
  .ZN(_038_)
);

AOI21_X1 _227_ (
  .A(_081_),
  .B1(_075_),
  .B2(_038_),
  .ZN(_039_)
);

AOI21_X1 _228_ (
  .A(_034_),
  .B1(_036_),
  .B2(_039_),
  .ZN(_008_)
);

NAND3_X1 _229_ (
  .A1(_028_),
  .A2(_065_),
  .A3(_108_),
  .ZN(_040_)
);

NAND3_X1 _230_ (
  .A1(_030_),
  .A2(_066_),
  .A3(_111_),
  .ZN(_041_)
);

NAND3_X1 _231_ (
  .A1(_040_),
  .A2(_041_),
  .A3(_079_),
  .ZN(_042_)
);

NAND2_X1 _232_ (
  .A1(_081_),
  .A2(\coef[30] ),
  .ZN(_043_)
);

NAND2_X1 _233_ (
  .A1(_042_),
  .A2(_043_),
  .ZN(_009_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_121_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_120_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_119_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_118_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_117_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_116_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_115_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_114_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_113_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_112_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$26ce9ce45d1136272d6a188b0b22329681d6199b\dctu

module \$paramod$16cad72ebc555f93621a2c70f423f14f85bbeb07\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _184_ (
  .A(x[1]),
  .ZN(_167_)
);

INV_X1 _185_ (
  .A(x[0]),
  .ZN(_166_)
);

BUF_X2 _186_ (
  .A(ena),
  .Z(_097_)
);

INV_X1 _187_ (
  .A(_097_),
  .ZN(_098_)
);

BUF_X2 _188_ (
  .A(y[2]),
  .Z(_099_)
);

INV_X2 _189_ (
  .A(_099_),
  .ZN(_100_)
);

INV_X2 _190_ (
  .A(x[2]),
  .ZN(_101_)
);

BUF_X8 _191_ (
  .A(_101_),
  .Z(_102_)
);

NAND2_X2 _192_ (
  .A1(_102_),
  .A2(_174_),
  .ZN(_103_)
);

INV_X1 _193_ (
  .A(_176_),
  .ZN(_104_)
);

BUF_X4 _194_ (
  .A(x[2]),
  .Z(_105_)
);

NAND2_X1 _195_ (
  .A1(_104_),
  .A2(_105_),
  .ZN(_106_)
);

BUF_X4 _196_ (
  .A(y[0]),
  .Z(_107_)
);

BUF_X4 _197_ (
  .A(_107_),
  .Z(_108_)
);

NAND3_X1 _198_ (
  .A1(_103_),
  .A2(_106_),
  .A3(_108_),
  .ZN(_109_)
);

INV_X1 _199_ (
  .A(y[0]),
  .ZN(_110_)
);

NAND2_X1 _200_ (
  .A1(_110_),
  .A2(_105_),
  .ZN(_111_)
);

BUF_X4 _201_ (
  .A(y[1]),
  .Z(_112_)
);

NAND2_X1 _202_ (
  .A1(_111_),
  .A2(_112_),
  .ZN(_113_)
);

INV_X1 _203_ (
  .A(_113_),
  .ZN(_114_)
);

AOI21_X1 _204_ (
  .A(_100_),
  .B1(_109_),
  .B2(_114_),
  .ZN(_115_)
);

INV_X1 _205_ (
  .A(_182_),
  .ZN(_116_)
);

NAND2_X2 _206_ (
  .A1(_102_),
  .A2(_116_),
  .ZN(_117_)
);

BUF_X4 _207_ (
  .A(_110_),
  .Z(_118_)
);

NAND2_X1 _208_ (
  .A1(_105_),
  .A2(_168_),
  .ZN(_119_)
);

NAND3_X2 _209_ (
  .A1(_117_),
  .A2(_118_),
  .A3(_119_),
  .ZN(_120_)
);

NAND2_X1 _210_ (
  .A1(_107_),
  .A2(x[0]),
  .ZN(_121_)
);

NAND2_X1 _211_ (
  .A1(_120_),
  .A2(_121_),
  .ZN(_122_)
);

INV_X4 _212_ (
  .A(_112_),
  .ZN(_123_)
);

BUF_X4 _213_ (
  .A(_123_),
  .Z(_124_)
);

NAND2_X1 _214_ (
  .A1(_122_),
  .A2(_124_),
  .ZN(_125_)
);

AOI21_X1 _215_ (
  .A(_098_),
  .B1(_115_),
  .B2(_125_),
  .ZN(_126_)
);

BUF_X4 _216_ (
  .A(_112_),
  .Z(_127_)
);

INV_X1 _217_ (
  .A(_172_),
  .ZN(_128_)
);

NAND2_X1 _218_ (
  .A1(_102_),
  .A2(_128_),
  .ZN(_129_)
);

NAND2_X1 _219_ (
  .A1(_105_),
  .A2(_178_),
  .ZN(_130_)
);

NAND3_X1 _220_ (
  .A1(_129_),
  .A2(_118_),
  .A3(_130_),
  .ZN(_131_)
);

NAND2_X1 _221_ (
  .A1(_101_),
  .A2(_107_),
  .ZN(_132_)
);

AOI21_X1 _222_ (
  .A(_127_),
  .B1(_131_),
  .B2(_132_),
  .ZN(_133_)
);

NAND2_X2 _223_ (
  .A1(_102_),
  .A2(_180_),
  .ZN(_134_)
);

INV_X1 _224_ (
  .A(_170_),
  .ZN(_135_)
);

NAND2_X1 _225_ (
  .A1(_135_),
  .A2(_105_),
  .ZN(_136_)
);

NAND3_X2 _226_ (
  .A1(_134_),
  .A2(_136_),
  .A3(_107_),
  .ZN(_137_)
);

AOI21_X1 _227_ (
  .A(_123_),
  .B1(_166_),
  .B2(_110_),
  .ZN(_138_)
);

NAND2_X1 _228_ (
  .A1(_137_),
  .A2(_138_),
  .ZN(_139_)
);

INV_X1 _229_ (
  .A(_139_),
  .ZN(_140_)
);

OAI21_X1 _230_ (
  .A(_100_),
  .B1(_133_),
  .B2(_140_),
  .ZN(_141_)
);

NAND2_X1 _231_ (
  .A1(_126_),
  .A2(_141_),
  .ZN(_142_)
);

NAND2_X1 _232_ (
  .A1(_098_),
  .A2(\coef[21] ),
  .ZN(_143_)
);

NAND2_X1 _233_ (
  .A1(_142_),
  .A2(_143_),
  .ZN(_000_)
);

NOR2_X1 _234_ (
  .A1(_097_),
  .A2(\coef[23] ),
  .ZN(_144_)
);

NAND2_X1 _235_ (
  .A1(_103_),
  .A2(_106_),
  .ZN(_145_)
);

NAND2_X1 _236_ (
  .A1(_145_),
  .A2(_118_),
  .ZN(_146_)
);

NAND2_X1 _237_ (
  .A1(_129_),
  .A2(_130_),
  .ZN(_147_)
);

NAND2_X2 _238_ (
  .A1(_147_),
  .A2(_108_),
  .ZN(_148_)
);

NAND3_X1 _239_ (
  .A1(_146_),
  .A2(_148_),
  .A3(_127_),
  .ZN(_149_)
);

NAND2_X1 _240_ (
  .A1(_111_),
  .A2(_121_),
  .ZN(_150_)
);

AOI21_X1 _241_ (
  .A(_100_),
  .B1(_150_),
  .B2(_124_),
  .ZN(_151_)
);

AOI21_X1 _242_ (
  .A(_098_),
  .B1(_149_),
  .B2(_151_),
  .ZN(_152_)
);

NAND3_X1 _243_ (
  .A1(_146_),
  .A2(_148_),
  .A3(_124_),
  .ZN(_153_)
);

OAI21_X1 _244_ (
  .A(_132_),
  .B1(_107_),
  .B2(x[0]),
  .ZN(_154_)
);

NAND2_X1 _245_ (
  .A1(_154_),
  .A2(_127_),
  .ZN(_155_)
);

NAND3_X1 _246_ (
  .A1(_153_),
  .A2(_100_),
  .A3(_155_),
  .ZN(_156_)
);

AOI21_X1 _247_ (
  .A(_144_),
  .B1(_152_),
  .B2(_156_),
  .ZN(_001_)
);

NOR2_X1 _248_ (
  .A1(_097_),
  .A2(\coef[24] ),
  .ZN(_009_)
);

AOI21_X1 _249_ (
  .A(_112_),
  .B1(_102_),
  .B2(_107_),
  .ZN(_010_)
);

AOI21_X1 _250_ (
  .A(_099_),
  .B1(_146_),
  .B2(_010_),
  .ZN(_011_)
);

XNOR2_X2 _251_ (
  .A(_105_),
  .B(_169_),
  .ZN(_012_)
);

NAND2_X1 _252_ (
  .A1(_012_),
  .A2(_108_),
  .ZN(_013_)
);

NAND2_X2 _253_ (
  .A1(_102_),
  .A2(_168_),
  .ZN(_014_)
);

NAND2_X1 _254_ (
  .A1(_116_),
  .A2(_105_),
  .ZN(_015_)
);

NAND3_X1 _255_ (
  .A1(_014_),
  .A2(_015_),
  .A3(_110_),
  .ZN(_016_)
);

NAND3_X1 _256_ (
  .A1(_013_),
  .A2(_127_),
  .A3(_016_),
  .ZN(_017_)
);

AOI21_X1 _257_ (
  .A(_098_),
  .B1(_011_),
  .B2(_017_),
  .ZN(_018_)
);

OR2_X4 _258_ (
  .A1(_012_),
  .A2(_108_),
  .ZN(_019_)
);

NAND2_X2 _259_ (
  .A1(_102_),
  .A2(_135_),
  .ZN(_020_)
);

NAND2_X1 _260_ (
  .A1(_105_),
  .A2(_180_),
  .ZN(_021_)
);

NAND3_X1 _261_ (
  .A1(_020_),
  .A2(_107_),
  .A3(_021_),
  .ZN(_022_)
);

NAND3_X1 _262_ (
  .A1(_019_),
  .A2(_124_),
  .A3(_022_),
  .ZN(_023_)
);

AOI21_X1 _263_ (
  .A(_100_),
  .B1(_148_),
  .B2(_114_),
  .ZN(_024_)
);

NAND2_X1 _264_ (
  .A1(_023_),
  .A2(_024_),
  .ZN(_025_)
);

AOI21_X2 _265_ (
  .A(_009_),
  .B1(_018_),
  .B2(_025_),
  .ZN(_002_)
);

NAND2_X1 _266_ (
  .A1(_120_),
  .A2(_022_),
  .ZN(_026_)
);

NAND2_X1 _267_ (
  .A1(_026_),
  .A2(_124_),
  .ZN(_027_)
);

NAND2_X1 _268_ (
  .A1(_102_),
  .A2(_178_),
  .ZN(_028_)
);

NAND2_X1 _269_ (
  .A1(_128_),
  .A2(_105_),
  .ZN(_029_)
);

NAND3_X1 _270_ (
  .A1(_028_),
  .A2(_029_),
  .A3(_108_),
  .ZN(_030_)
);

NAND3_X1 _271_ (
  .A1(_030_),
  .A2(_131_),
  .A3(_127_),
  .ZN(_031_)
);

NAND3_X1 _272_ (
  .A1(_027_),
  .A2(_031_),
  .A3(_100_),
  .ZN(_032_)
);

NAND2_X1 _273_ (
  .A1(_137_),
  .A2(_016_),
  .ZN(_033_)
);

NAND2_X1 _274_ (
  .A1(_033_),
  .A2(_127_),
  .ZN(_034_)
);

NAND2_X1 _275_ (
  .A1(_102_),
  .A2(_104_),
  .ZN(_035_)
);

NAND2_X1 _276_ (
  .A1(_105_),
  .A2(_174_),
  .ZN(_036_)
);

NAND3_X1 _277_ (
  .A1(_035_),
  .A2(_118_),
  .A3(_036_),
  .ZN(_037_)
);

NAND3_X1 _278_ (
  .A1(_109_),
  .A2(_037_),
  .A3(_124_),
  .ZN(_038_)
);

NAND3_X1 _279_ (
  .A1(_034_),
  .A2(_038_),
  .A3(_099_),
  .ZN(_039_)
);

NAND3_X1 _280_ (
  .A1(_032_),
  .A2(_039_),
  .A3(_097_),
  .ZN(_040_)
);

NAND2_X1 _281_ (
  .A1(_098_),
  .A2(\coef[10] ),
  .ZN(_041_)
);

NAND2_X1 _282_ (
  .A1(_040_),
  .A2(_041_),
  .ZN(_003_)
);

NOR2_X1 _283_ (
  .A1(_097_),
  .A2(\coef[26] ),
  .ZN(_042_)
);

NAND2_X1 _284_ (
  .A1(_166_),
  .A2(_107_),
  .ZN(_043_)
);

OAI21_X1 _285_ (
  .A(_100_),
  .B1(_043_),
  .B2(_112_),
  .ZN(_044_)
);

NOR2_X1 _286_ (
  .A1(_108_),
  .A2(_112_),
  .ZN(_045_)
);

NAND2_X1 _287_ (
  .A1(_134_),
  .A2(_136_),
  .ZN(_046_)
);

AOI21_X1 _288_ (
  .A(_044_),
  .B1(_045_),
  .B2(_046_),
  .ZN(_047_)
);

NAND3_X1 _289_ (
  .A1(_146_),
  .A2(_127_),
  .A3(_043_),
  .ZN(_048_)
);

AOI21_X1 _290_ (
  .A(_098_),
  .B1(_047_),
  .B2(_048_),
  .ZN(_049_)
);

NAND3_X1 _291_ (
  .A1(_117_),
  .A2(_108_),
  .A3(_119_),
  .ZN(_050_)
);

AOI21_X1 _292_ (
  .A(_100_),
  .B1(_050_),
  .B2(_138_),
  .ZN(_051_)
);

OAI21_X1 _293_ (
  .A(_148_),
  .B1(_108_),
  .B2(_166_),
  .ZN(_052_)
);

OAI21_X1 _294_ (
  .A(_051_),
  .B1(_052_),
  .B2(_127_),
  .ZN(_053_)
);

AOI21_X2 _295_ (
  .A(_042_),
  .B1(_049_),
  .B2(_053_),
  .ZN(_004_)
);

NOR2_X1 _296_ (
  .A1(_097_),
  .A2(\coef[13] ),
  .ZN(_054_)
);

NAND2_X1 _297_ (
  .A1(_028_),
  .A2(_029_),
  .ZN(_055_)
);

NAND2_X1 _298_ (
  .A1(_055_),
  .A2(_118_),
  .ZN(_056_)
);

NAND3_X1 _299_ (
  .A1(_013_),
  .A2(_056_),
  .A3(_124_),
  .ZN(_057_)
);

NOR2_X1 _300_ (
  .A1(_107_),
  .A2(x[1]),
  .ZN(_058_)
);

NOR2_X1 _301_ (
  .A1(_058_),
  .A2(_123_),
  .ZN(_059_)
);

AOI21_X1 _302_ (
  .A(_100_),
  .B1(_022_),
  .B2(_059_),
  .ZN(_060_)
);

AOI21_X1 _303_ (
  .A(_098_),
  .B1(_057_),
  .B2(_060_),
  .ZN(_061_)
);

NAND2_X1 _304_ (
  .A1(_107_),
  .A2(x[1]),
  .ZN(_062_)
);

NAND2_X1 _305_ (
  .A1(_062_),
  .A2(_124_),
  .ZN(_063_)
);

INV_X1 _306_ (
  .A(_063_),
  .ZN(_064_)
);

AOI21_X1 _307_ (
  .A(_099_),
  .B1(_016_),
  .B2(_064_),
  .ZN(_065_)
);

NAND2_X1 _308_ (
  .A1(_019_),
  .A2(_127_),
  .ZN(_066_)
);

AOI21_X1 _309_ (
  .A(_118_),
  .B1(_035_),
  .B2(_036_),
  .ZN(_067_)
);

OAI21_X1 _310_ (
  .A(_065_),
  .B1(_066_),
  .B2(_067_),
  .ZN(_068_)
);

AOI21_X2 _311_ (
  .A(_054_),
  .B1(_061_),
  .B2(_068_),
  .ZN(_005_)
);

OAI21_X1 _312_ (
  .A(_099_),
  .B1(_150_),
  .B2(_123_),
  .ZN(_069_)
);

INV_X1 _313_ (
  .A(_069_),
  .ZN(_070_)
);

INV_X1 _314_ (
  .A(_062_),
  .ZN(_071_)
);

AOI21_X1 _315_ (
  .A(_071_),
  .B1(_012_),
  .B2(_118_),
  .ZN(_072_)
);

OAI21_X1 _316_ (
  .A(_070_),
  .B1(_072_),
  .B2(_127_),
  .ZN(_073_)
);

OAI21_X1 _317_ (
  .A(_059_),
  .B1(_012_),
  .B2(_118_),
  .ZN(_074_)
);

NAND2_X1 _318_ (
  .A1(_154_),
  .A2(_124_),
  .ZN(_075_)
);

NAND2_X1 _319_ (
  .A1(_074_),
  .A2(_075_),
  .ZN(_076_)
);

NAND2_X1 _320_ (
  .A1(_076_),
  .A2(_100_),
  .ZN(_077_)
);

NAND2_X1 _321_ (
  .A1(_073_),
  .A2(_077_),
  .ZN(_078_)
);

NAND2_X2 _322_ (
  .A1(_078_),
  .A2(_097_),
  .ZN(_079_)
);

NAND2_X1 _323_ (
  .A1(_098_),
  .A2(\coef[28] ),
  .ZN(_080_)
);

NAND2_X2 _324_ (
  .A1(_079_),
  .A2(_080_),
  .ZN(_006_)
);

NAND3_X1 _325_ (
  .A1(_020_),
  .A2(_118_),
  .A3(_021_),
  .ZN(_081_)
);

NAND3_X1 _326_ (
  .A1(_137_),
  .A2(_081_),
  .A3(_124_),
  .ZN(_082_)
);

NAND2_X1 _327_ (
  .A1(_114_),
  .A2(_062_),
  .ZN(_083_)
);

NAND3_X1 _328_ (
  .A1(_082_),
  .A2(_099_),
  .A3(_083_),
  .ZN(_084_)
);

NAND3_X1 _329_ (
  .A1(_014_),
  .A2(_015_),
  .A3(_108_),
  .ZN(_085_)
);

NAND3_X1 _330_ (
  .A1(_085_),
  .A2(_120_),
  .A3(_112_),
  .ZN(_086_)
);

INV_X1 _331_ (
  .A(_058_),
  .ZN(_087_)
);

AOI21_X1 _332_ (
  .A(_099_),
  .B1(_010_),
  .B2(_087_),
  .ZN(_088_)
);

NAND2_X1 _333_ (
  .A1(_086_),
  .A2(_088_),
  .ZN(_089_)
);

NAND2_X1 _334_ (
  .A1(_084_),
  .A2(_089_),
  .ZN(_090_)
);

NAND2_X1 _335_ (
  .A1(_090_),
  .A2(_097_),
  .ZN(_091_)
);

NAND2_X1 _336_ (
  .A1(_098_),
  .A2(\coef[29] ),
  .ZN(_092_)
);

NAND2_X1 _337_ (
  .A1(_091_),
  .A2(_092_),
  .ZN(_007_)
);

NOR2_X1 _338_ (
  .A1(_097_),
  .A2(\coef[30] ),
  .ZN(_093_)
);

OAI21_X1 _339_ (
  .A(_099_),
  .B1(_118_),
  .B2(_123_),
  .ZN(_094_)
);

OAI21_X1 _340_ (
  .A(_094_),
  .B1(_108_),
  .B2(_112_),
  .ZN(_095_)
);

XNOR2_X1 _341_ (
  .A(_095_),
  .B(_102_),
  .ZN(_096_)
);

AOI21_X1 _342_ (
  .A(_093_),
  .B1(_096_),
  .B2(_097_),
  .ZN(_008_)
);

HA_X1 _343_ (
  .A(_166_),
  .B(_167_),
  .CO(_168_),
  .S(_169_)
);

HA_X1 _344_ (
  .A(_166_),
  .B(_167_),
  .CO(_170_),
  .S(_171_)
);

HA_X1 _345_ (
  .A(_166_),
  .B(x[1]),
  .CO(_172_),
  .S(_173_)
);

HA_X1 _346_ (
  .A(_166_),
  .B(x[1]),
  .CO(_174_),
  .S(_175_)
);

HA_X1 _347_ (
  .A(x[0]),
  .B(_167_),
  .CO(_176_),
  .S(_177_)
);

HA_X1 _348_ (
  .A(x[0]),
  .B(_167_),
  .CO(_178_),
  .S(_179_)
);

HA_X1 _349_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_180_),
  .S(_181_)
);

HA_X1 _350_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_182_),
  .S(_183_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_165_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_164_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_163_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_162_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_161_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_160_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_159_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_158_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_157_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$16cad72ebc555f93621a2c70f423f14f85bbeb07\dctu

module \$paramod$022e4835c44d221125856d68f8603b7186431212\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire \coef[10] ;
wire \coef[11] ;
wire \coef[13] ;
wire \coef[15] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

BUF_X4 _30_ (
  .A(x[2]),
  .Z(_04_)
);

INV_X4 _31_ (
  .A(_04_),
  .ZN(_05_)
);

INV_X1 _32_ (
  .A(x[0]),
  .ZN(_06_)
);

NAND2_X1 _33_ (
  .A1(_05_),
  .A2(_06_),
  .ZN(_07_)
);

BUF_X4 _34_ (
  .A(ena),
  .Z(_08_)
);

NAND2_X1 _35_ (
  .A1(_04_),
  .A2(x[0]),
  .ZN(_09_)
);

NAND3_X1 _36_ (
  .A1(_07_),
  .A2(_08_),
  .A3(_09_),
  .ZN(_10_)
);

INV_X1 _37_ (
  .A(_08_),
  .ZN(_11_)
);

NAND2_X1 _38_ (
  .A1(_11_),
  .A2(\coef[13] ),
  .ZN(_12_)
);

NAND2_X1 _39_ (
  .A1(_10_),
  .A2(_12_),
  .ZN(_00_)
);

INV_X1 _40_ (
  .A(x[1]),
  .ZN(_13_)
);

NAND2_X1 _41_ (
  .A1(_05_),
  .A2(_13_),
  .ZN(_14_)
);

NAND2_X1 _42_ (
  .A1(_04_),
  .A2(x[1]),
  .ZN(_15_)
);

NAND3_X1 _43_ (
  .A1(_14_),
  .A2(_08_),
  .A3(_15_),
  .ZN(_16_)
);

NAND2_X1 _44_ (
  .A1(_11_),
  .A2(\coef[15] ),
  .ZN(_17_)
);

NAND2_X1 _45_ (
  .A1(_16_),
  .A2(_17_),
  .ZN(_01_)
);

NAND2_X1 _46_ (
  .A1(_06_),
  .A2(_04_),
  .ZN(_18_)
);

NAND2_X2 _47_ (
  .A1(_05_),
  .A2(x[0]),
  .ZN(_19_)
);

NAND3_X1 _48_ (
  .A1(_18_),
  .A2(_19_),
  .A3(_08_),
  .ZN(_20_)
);

NAND2_X1 _49_ (
  .A1(_11_),
  .A2(\coef[10] ),
  .ZN(_21_)
);

NAND2_X1 _50_ (
  .A1(_20_),
  .A2(_21_),
  .ZN(_02_)
);

NAND2_X1 _51_ (
  .A1(_13_),
  .A2(_04_),
  .ZN(_22_)
);

NAND2_X2 _52_ (
  .A1(_05_),
  .A2(x[1]),
  .ZN(_23_)
);

NAND3_X1 _53_ (
  .A1(_22_),
  .A2(_23_),
  .A3(_08_),
  .ZN(_24_)
);

NAND2_X1 _54_ (
  .A1(_11_),
  .A2(\coef[11] ),
  .ZN(_25_)
);

NAND2_X1 _55_ (
  .A1(_24_),
  .A2(_25_),
  .ZN(_03_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_03_),
  .CK(clk),
  .Q(\coef[11] ),
  .QN(_26_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_29_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_02_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_27_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_01_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_28_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[15] , \coef[15] , \coef[10] , \coef[13] , \coef[10] , \coef[15] , \coef[15] , \coef[11] , \coef[10] , \coef[11] , \coef[15] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$022e4835c44d221125856d68f8603b7186431212\dctu

module \$paramod$141b5017b00a41bd6bcdd772ef8ad836aaf4019f\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _070_ (
  .A(x[1]),
  .ZN(_008_)
);

INV_X2 _071_ (
  .A(x[0]),
  .ZN(_009_)
);

NAND2_X2 _072_ (
  .A1(_008_),
  .A2(_009_),
  .ZN(_010_)
);

NAND2_X1 _073_ (
  .A1(x[1]),
  .A2(x[0]),
  .ZN(_011_)
);

NAND2_X2 _074_ (
  .A1(_010_),
  .A2(_011_),
  .ZN(_012_)
);

BUF_X1 _075_ (
  .A(y[1]),
  .Z(_013_)
);

NAND2_X1 _076_ (
  .A1(_012_),
  .A2(_013_),
  .ZN(_014_)
);

NAND2_X1 _077_ (
  .A1(_008_),
  .A2(x[0]),
  .ZN(_015_)
);

NAND2_X1 _078_ (
  .A1(_009_),
  .A2(x[1]),
  .ZN(_016_)
);

NAND2_X2 _079_ (
  .A1(_015_),
  .A2(_016_),
  .ZN(_017_)
);

INV_X1 _080_ (
  .A(_013_),
  .ZN(_018_)
);

NAND2_X1 _081_ (
  .A1(_017_),
  .A2(_018_),
  .ZN(_019_)
);

CLKBUF_X3 _082_ (
  .A(ena),
  .Z(_020_)
);

NAND3_X1 _083_ (
  .A1(_014_),
  .A2(_019_),
  .A3(_020_),
  .ZN(_021_)
);

INV_X1 _084_ (
  .A(\coef[21] ),
  .ZN(_022_)
);

OAI21_X1 _085_ (
  .A(_021_),
  .B1(_022_),
  .B2(_020_),
  .ZN(_000_)
);

NAND2_X2 _086_ (
  .A1(_012_),
  .A2(y[0]),
  .ZN(_023_)
);

INV_X1 _087_ (
  .A(y[0]),
  .ZN(_024_)
);

NAND3_X1 _088_ (
  .A1(_010_),
  .A2(_024_),
  .A3(_011_),
  .ZN(_025_)
);

NAND3_X2 _089_ (
  .A1(_023_),
  .A2(_025_),
  .A3(_013_),
  .ZN(_026_)
);

CLKBUF_X3 _090_ (
  .A(y[2]),
  .Z(_027_)
);

INV_X1 _091_ (
  .A(_027_),
  .ZN(_028_)
);

NAND2_X1 _092_ (
  .A1(_012_),
  .A2(_018_),
  .ZN(_029_)
);

NAND3_X2 _093_ (
  .A1(_026_),
  .A2(_028_),
  .A3(_029_),
  .ZN(_030_)
);

NAND3_X2 _094_ (
  .A1(_023_),
  .A2(_025_),
  .A3(_018_),
  .ZN(_031_)
);

NAND2_X1 _095_ (
  .A1(_017_),
  .A2(_013_),
  .ZN(_032_)
);

NAND3_X2 _096_ (
  .A1(_031_),
  .A2(_027_),
  .A3(_032_),
  .ZN(_033_)
);

NAND2_X1 _097_ (
  .A1(_030_),
  .A2(_033_),
  .ZN(_034_)
);

NAND2_X1 _098_ (
  .A1(_034_),
  .A2(_020_),
  .ZN(_035_)
);

INV_X1 _099_ (
  .A(ena),
  .ZN(_036_)
);

NAND2_X1 _100_ (
  .A1(_036_),
  .A2(\coef[22] ),
  .ZN(_037_)
);

NAND2_X2 _101_ (
  .A1(_035_),
  .A2(_037_),
  .ZN(_001_)
);

NAND3_X1 _102_ (
  .A1(_026_),
  .A2(_027_),
  .A3(_019_),
  .ZN(_038_)
);

NAND3_X1 _103_ (
  .A1(_031_),
  .A2(_028_),
  .A3(_014_),
  .ZN(_039_)
);

NAND3_X1 _104_ (
  .A1(_038_),
  .A2(_039_),
  .A3(_020_),
  .ZN(_040_)
);

NAND2_X1 _105_ (
  .A1(_036_),
  .A2(\coef[23] ),
  .ZN(_041_)
);

NAND2_X1 _106_ (
  .A1(_040_),
  .A2(_041_),
  .ZN(_002_)
);

NAND3_X1 _107_ (
  .A1(_030_),
  .A2(_033_),
  .A3(_020_),
  .ZN(_042_)
);

NAND2_X1 _108_ (
  .A1(_036_),
  .A2(\coef[14] ),
  .ZN(_043_)
);

NAND2_X1 _109_ (
  .A1(_042_),
  .A2(_043_),
  .ZN(_003_)
);

NOR2_X1 _110_ (
  .A1(_020_),
  .A2(\coef[13] ),
  .ZN(_044_)
);

XNOR2_X1 _111_ (
  .A(_017_),
  .B(_027_),
  .ZN(_045_)
);

AOI21_X1 _112_ (
  .A(_044_),
  .B1(_045_),
  .B2(_020_),
  .ZN(_004_)
);

NAND2_X2 _113_ (
  .A1(_017_),
  .A2(y[0]),
  .ZN(_046_)
);

NAND2_X2 _114_ (
  .A1(_012_),
  .A2(_024_),
  .ZN(_047_)
);

NAND3_X1 _115_ (
  .A1(_046_),
  .A2(_047_),
  .A3(_013_),
  .ZN(_048_)
);

NAND3_X1 _116_ (
  .A1(_048_),
  .A2(_031_),
  .A3(_027_),
  .ZN(_049_)
);

NAND3_X1 _117_ (
  .A1(_046_),
  .A2(_047_),
  .A3(_018_),
  .ZN(_050_)
);

NAND3_X1 _118_ (
  .A1(_050_),
  .A2(_026_),
  .A3(_028_),
  .ZN(_051_)
);

NAND3_X1 _119_ (
  .A1(_049_),
  .A2(_051_),
  .A3(_020_),
  .ZN(_052_)
);

NAND2_X1 _120_ (
  .A1(_036_),
  .A2(\coef[28] ),
  .ZN(_053_)
);

NAND2_X1 _121_ (
  .A1(_052_),
  .A2(_053_),
  .ZN(_005_)
);

NAND3_X1 _122_ (
  .A1(_050_),
  .A2(_027_),
  .A3(_032_),
  .ZN(_054_)
);

NAND3_X1 _123_ (
  .A1(_048_),
  .A2(_028_),
  .A3(_029_),
  .ZN(_055_)
);

NAND3_X1 _124_ (
  .A1(_054_),
  .A2(_055_),
  .A3(_020_),
  .ZN(_056_)
);

NAND2_X1 _125_ (
  .A1(_036_),
  .A2(\coef[15] ),
  .ZN(_057_)
);

NAND2_X1 _126_ (
  .A1(_056_),
  .A2(_057_),
  .ZN(_006_)
);

NAND3_X1 _127_ (
  .A1(_048_),
  .A2(_027_),
  .A3(_019_),
  .ZN(_058_)
);

NAND3_X1 _128_ (
  .A1(_050_),
  .A2(_028_),
  .A3(_014_),
  .ZN(_059_)
);

NAND3_X1 _129_ (
  .A1(_058_),
  .A2(_059_),
  .A3(_020_),
  .ZN(_060_)
);

NAND2_X1 _130_ (
  .A1(_036_),
  .A2(\coef[12] ),
  .ZN(_061_)
);

NAND2_X1 _131_ (
  .A1(_060_),
  .A2(_061_),
  .ZN(_007_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_069_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_068_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_067_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_066_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_065_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_064_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_063_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_062_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$141b5017b00a41bd6bcdd772ef8ad836aaf4019f\dctu

module \$paramod$2ce29d501700894abc3f54c094daafc2d8c2c211\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire \coef[10] ;
wire \coef[11] ;
wire \coef[13] ;
wire \coef[15] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

NOR2_X1 _33_ (
  .A1(\coef[11] ),
  .A2(ena),
  .ZN(_04_)
);

INV_X1 _34_ (
  .A(ena),
  .ZN(_05_)
);

INV_X1 _35_ (
  .A(x[1]),
  .ZN(_06_)
);

INV_X1 _36_ (
  .A(x[0]),
  .ZN(_07_)
);

NAND2_X2 _37_ (
  .A1(_06_),
  .A2(_07_),
  .ZN(_08_)
);

NAND2_X1 _38_ (
  .A1(x[1]),
  .A2(x[0]),
  .ZN(_09_)
);

NAND2_X4 _39_ (
  .A1(_08_),
  .A2(_09_),
  .ZN(_10_)
);

INV_X1 _40_ (
  .A(y[0]),
  .ZN(_11_)
);

INV_X2 _41_ (
  .A(y[2]),
  .ZN(_12_)
);

NAND2_X4 _42_ (
  .A1(_11_),
  .A2(_12_),
  .ZN(_13_)
);

NAND2_X1 _43_ (
  .A1(y[0]),
  .A2(y[2]),
  .ZN(_14_)
);

NAND2_X4 _44_ (
  .A1(_13_),
  .A2(_14_),
  .ZN(_15_)
);

AOI21_X4 _45_ (
  .A(_05_),
  .B1(_10_),
  .B2(_15_),
  .ZN(_16_)
);

OR2_X4 _46_ (
  .A1(_15_),
  .A2(_10_),
  .ZN(_17_)
);

AOI21_X4 _47_ (
  .A(_04_),
  .B1(_16_),
  .B2(_17_),
  .ZN(_00_)
);

NOR2_X1 _48_ (
  .A1(ena),
  .A2(\coef[13] ),
  .ZN(_18_)
);

INV_X1 _49_ (
  .A(y[1]),
  .ZN(_19_)
);

NAND2_X2 _50_ (
  .A1(_12_),
  .A2(_19_),
  .ZN(_20_)
);

NAND2_X1 _51_ (
  .A1(y[2]),
  .A2(y[1]),
  .ZN(_21_)
);

NAND2_X2 _52_ (
  .A1(_20_),
  .A2(_21_),
  .ZN(_22_)
);

AOI21_X2 _53_ (
  .A(_05_),
  .B1(_10_),
  .B2(_22_),
  .ZN(_23_)
);

OR2_X4 _54_ (
  .A1(_22_),
  .A2(_10_),
  .ZN(_24_)
);

AOI21_X2 _55_ (
  .A(_18_),
  .B1(_23_),
  .B2(_24_),
  .ZN(_01_)
);

NAND2_X2 _56_ (
  .A1(_23_),
  .A2(_24_),
  .ZN(_25_)
);

NAND2_X1 _57_ (
  .A1(_05_),
  .A2(\coef[10] ),
  .ZN(_26_)
);

NAND2_X2 _58_ (
  .A1(_25_),
  .A2(_26_),
  .ZN(_02_)
);

NAND2_X4 _59_ (
  .A1(_16_),
  .A2(_17_),
  .ZN(_27_)
);

NAND2_X1 _60_ (
  .A1(_05_),
  .A2(\coef[15] ),
  .ZN(_28_)
);

NAND2_X2 _61_ (
  .A1(_27_),
  .A2(_28_),
  .ZN(_03_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[11] ),
  .QN(_32_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_01_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_31_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_02_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_30_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_03_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_29_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[15] , \coef[15] , \coef[10] , \coef[13] , \coef[10] , \coef[15] , \coef[15] , \coef[11] , \coef[10] , \coef[11] , \coef[15] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$2ce29d501700894abc3f54c094daafc2d8c2c211\dctu

module \$paramod$30e2d72cbb2d6c7d2f48769e891fec5593e1f756\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _057_ (
  .A(x[0]),
  .ZN(_047_)
);

INV_X1 _058_ (
  .A(x[1]),
  .ZN(_048_)
);

INV_X1 _059_ (
  .A(_051_),
  .ZN(_008_)
);

BUF_X4 _060_ (
  .A(x[2]),
  .Z(_009_)
);

NAND2_X1 _061_ (
  .A1(_008_),
  .A2(_009_),
  .ZN(_010_)
);

INV_X4 _062_ (
  .A(_009_),
  .ZN(_011_)
);

NAND2_X1 _063_ (
  .A1(_011_),
  .A2(_053_),
  .ZN(_012_)
);

BUF_X4 _064_ (
  .A(ena),
  .Z(_013_)
);

NAND3_X1 _065_ (
  .A1(_010_),
  .A2(_012_),
  .A3(_013_),
  .ZN(_014_)
);

INV_X4 _066_ (
  .A(_013_),
  .ZN(_015_)
);

BUF_X16 _067_ (
  .A(_015_),
  .Z(_016_)
);

NAND2_X1 _068_ (
  .A1(_016_),
  .A2(\coef[13] ),
  .ZN(_017_)
);

NAND2_X1 _069_ (
  .A1(_014_),
  .A2(_017_),
  .ZN(_000_)
);

INV_X1 _070_ (
  .A(_050_),
  .ZN(_018_)
);

NAND2_X1 _071_ (
  .A1(_011_),
  .A2(_018_),
  .ZN(_019_)
);

NAND2_X1 _072_ (
  .A1(_009_),
  .A2(_050_),
  .ZN(_020_)
);

NAND3_X1 _073_ (
  .A1(_019_),
  .A2(_013_),
  .A3(_020_),
  .ZN(_021_)
);

NAND2_X1 _074_ (
  .A1(_016_),
  .A2(\coef[14] ),
  .ZN(_022_)
);

NAND2_X1 _075_ (
  .A1(_021_),
  .A2(_022_),
  .ZN(_001_)
);

NAND2_X2 _076_ (
  .A1(_016_),
  .A2(\coef[15] ),
  .ZN(_023_)
);

OAI21_X2 _077_ (
  .A(_023_),
  .B1(x[1]),
  .B2(_016_),
  .ZN(_002_)
);

NAND2_X2 _078_ (
  .A1(_016_),
  .A2(\coef[12] ),
  .ZN(_024_)
);

OAI21_X2 _079_ (
  .A(_024_),
  .B1(_011_),
  .B2(_016_),
  .ZN(_003_)
);

INV_X1 _080_ (
  .A(_049_),
  .ZN(_025_)
);

NAND2_X1 _081_ (
  .A1(_025_),
  .A2(_009_),
  .ZN(_026_)
);

NAND2_X1 _082_ (
  .A1(_011_),
  .A2(_055_),
  .ZN(_027_)
);

NAND3_X1 _083_ (
  .A1(_026_),
  .A2(_027_),
  .A3(_013_),
  .ZN(_028_)
);

NAND2_X1 _084_ (
  .A1(_016_),
  .A2(\coef[21] ),
  .ZN(_029_)
);

NAND2_X1 _085_ (
  .A1(_028_),
  .A2(_029_),
  .ZN(_004_)
);

NAND2_X1 _086_ (
  .A1(_018_),
  .A2(_009_),
  .ZN(_030_)
);

NAND2_X1 _087_ (
  .A1(_011_),
  .A2(_050_),
  .ZN(_031_)
);

NAND3_X1 _088_ (
  .A1(_030_),
  .A2(_031_),
  .A3(_013_),
  .ZN(_032_)
);

NAND2_X1 _089_ (
  .A1(_016_),
  .A2(\coef[22] ),
  .ZN(_033_)
);

NAND2_X1 _090_ (
  .A1(_032_),
  .A2(_033_),
  .ZN(_005_)
);

NAND2_X2 _091_ (
  .A1(_016_),
  .A2(\coef[23] ),
  .ZN(_034_)
);

OAI21_X2 _092_ (
  .A(_034_),
  .B1(_047_),
  .B2(_016_),
  .ZN(_006_)
);

NAND2_X1 _093_ (
  .A1(_015_),
  .A2(\coef[28] ),
  .ZN(_035_)
);

NAND2_X1 _094_ (
  .A1(_009_),
  .A2(_053_),
  .ZN(_036_)
);

NAND2_X1 _095_ (
  .A1(_036_),
  .A2(_013_),
  .ZN(_037_)
);

NOR2_X1 _096_ (
  .A1(_009_),
  .A2(_051_),
  .ZN(_038_)
);

OAI21_X1 _097_ (
  .A(_035_),
  .B1(_037_),
  .B2(_038_),
  .ZN(_007_)
);

HA_X1 _098_ (
  .A(_047_),
  .B(_048_),
  .CO(_049_),
  .S(_050_)
);

HA_X1 _099_ (
  .A(_047_),
  .B(x[1]),
  .CO(_051_),
  .S(_052_)
);

HA_X1 _100_ (
  .A(x[0]),
  .B(_048_),
  .CO(_053_),
  .S(_054_)
);

HA_X1 _101_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_055_),
  .S(_056_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_042_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_041_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_040_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_045_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_046_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_039_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_044_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_043_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$30e2d72cbb2d6c7d2f48769e891fec5593e1f756\dctu

module \$paramod$32a02d514417e24bb09b7885b9c053483ac7784d\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

BUF_X1 _103_ (
  .A(ena),
  .Z(_027_)
);

BUF_X1 _104_ (
  .A(_027_),
  .Z(_028_)
);

NOR2_X1 _105_ (
  .A1(\coef[15] ),
  .A2(_028_),
  .ZN(_029_)
);

INV_X1 _106_ (
  .A(_027_),
  .ZN(_030_)
);

INV_X2 _107_ (
  .A(x[2]),
  .ZN(_031_)
);

INV_X1 _108_ (
  .A(x[0]),
  .ZN(_032_)
);

NAND2_X4 _109_ (
  .A1(_031_),
  .A2(_032_),
  .ZN(_033_)
);

NAND2_X2 _110_ (
  .A1(x[2]),
  .A2(x[0]),
  .ZN(_034_)
);

NAND2_X4 _111_ (
  .A1(_033_),
  .A2(_034_),
  .ZN(_035_)
);

BUF_X2 _112_ (
  .A(y[1]),
  .Z(_036_)
);

INV_X2 _113_ (
  .A(_036_),
  .ZN(_037_)
);

NAND2_X1 _114_ (
  .A1(_035_),
  .A2(_037_),
  .ZN(_038_)
);

INV_X1 _115_ (
  .A(x[1]),
  .ZN(_039_)
);

NAND2_X2 _116_ (
  .A1(_031_),
  .A2(_039_),
  .ZN(_040_)
);

NAND2_X1 _117_ (
  .A1(x[2]),
  .A2(x[1]),
  .ZN(_041_)
);

NAND3_X1 _118_ (
  .A1(_040_),
  .A2(_036_),
  .A3(_041_),
  .ZN(_042_)
);

NAND2_X1 _119_ (
  .A1(_038_),
  .A2(_042_),
  .ZN(_043_)
);

BUF_X2 _120_ (
  .A(y[0]),
  .Z(_044_)
);

NAND2_X1 _121_ (
  .A1(_043_),
  .A2(_044_),
  .ZN(_045_)
);

INV_X2 _122_ (
  .A(_044_),
  .ZN(_046_)
);

NAND3_X2 _123_ (
  .A1(_033_),
  .A2(_046_),
  .A3(_034_),
  .ZN(_047_)
);

BUF_X1 _124_ (
  .A(y[2]),
  .Z(_048_)
);

AND2_X1 _125_ (
  .A1(_047_),
  .A2(_048_),
  .ZN(_049_)
);

AOI21_X1 _126_ (
  .A(_030_),
  .B1(_045_),
  .B2(_049_),
  .ZN(_050_)
);

NAND3_X2 _127_ (
  .A1(_040_),
  .A2(_046_),
  .A3(_041_),
  .ZN(_051_)
);

NAND3_X1 _128_ (
  .A1(_033_),
  .A2(_044_),
  .A3(_034_),
  .ZN(_052_)
);

NAND2_X1 _129_ (
  .A1(_051_),
  .A2(_052_),
  .ZN(_053_)
);

NAND2_X1 _130_ (
  .A1(_053_),
  .A2(_037_),
  .ZN(_054_)
);

NAND2_X2 _131_ (
  .A1(_035_),
  .A2(_044_),
  .ZN(_055_)
);

NAND3_X2 _132_ (
  .A1(_055_),
  .A2(_047_),
  .A3(_036_),
  .ZN(_056_)
);

NAND2_X1 _133_ (
  .A1(_054_),
  .A2(_056_),
  .ZN(_057_)
);

INV_X2 _134_ (
  .A(_048_),
  .ZN(_058_)
);

NAND2_X1 _135_ (
  .A1(_057_),
  .A2(_058_),
  .ZN(_059_)
);

AOI21_X2 _136_ (
  .A(_029_),
  .B1(_050_),
  .B2(_059_),
  .ZN(_000_)
);

NAND2_X1 _137_ (
  .A1(_039_),
  .A2(x[2]),
  .ZN(_060_)
);

NAND2_X2 _138_ (
  .A1(_031_),
  .A2(x[1]),
  .ZN(_061_)
);

NAND3_X2 _139_ (
  .A1(_060_),
  .A2(_061_),
  .A3(_044_),
  .ZN(_062_)
);

NAND2_X2 _140_ (
  .A1(_062_),
  .A2(_051_),
  .ZN(_063_)
);

NAND2_X2 _141_ (
  .A1(_063_),
  .A2(_036_),
  .ZN(_064_)
);

NAND3_X1 _142_ (
  .A1(_055_),
  .A2(_047_),
  .A3(_037_),
  .ZN(_065_)
);

NAND3_X1 _143_ (
  .A1(_064_),
  .A2(_065_),
  .A3(_048_),
  .ZN(_066_)
);

NAND3_X1 _144_ (
  .A1(_060_),
  .A2(_061_),
  .A3(_046_),
  .ZN(_067_)
);

NAND3_X1 _145_ (
  .A1(_040_),
  .A2(_044_),
  .A3(_041_),
  .ZN(_068_)
);

NAND3_X1 _146_ (
  .A1(_067_),
  .A2(_068_),
  .A3(_037_),
  .ZN(_069_)
);

NAND3_X1 _147_ (
  .A1(_056_),
  .A2(_069_),
  .A3(_058_),
  .ZN(_070_)
);

NAND3_X1 _148_ (
  .A1(_066_),
  .A2(_070_),
  .A3(_028_),
  .ZN(_071_)
);

NAND2_X1 _149_ (
  .A1(_030_),
  .A2(\coef[21] ),
  .ZN(_072_)
);

NAND2_X1 _150_ (
  .A1(_071_),
  .A2(_072_),
  .ZN(_001_)
);

NOR2_X1 _151_ (
  .A1(_028_),
  .A2(\coef[22] ),
  .ZN(_073_)
);

XNOR2_X1 _152_ (
  .A(_035_),
  .B(_058_),
  .ZN(_074_)
);

AOI21_X1 _153_ (
  .A(_073_),
  .B1(_074_),
  .B2(_028_),
  .ZN(_002_)
);

NAND3_X1 _154_ (
  .A1(_047_),
  .A2(_068_),
  .A3(_037_),
  .ZN(_075_)
);

NAND3_X1 _155_ (
  .A1(_062_),
  .A2(_051_),
  .A3(_036_),
  .ZN(_076_)
);

NAND3_X1 _156_ (
  .A1(_075_),
  .A2(_076_),
  .A3(_048_),
  .ZN(_077_)
);

NAND2_X1 _157_ (
  .A1(_053_),
  .A2(_036_),
  .ZN(_078_)
);

NAND3_X1 _158_ (
  .A1(_062_),
  .A2(_051_),
  .A3(_037_),
  .ZN(_079_)
);

NAND3_X1 _159_ (
  .A1(_078_),
  .A2(_079_),
  .A3(_058_),
  .ZN(_080_)
);

NAND3_X1 _160_ (
  .A1(_077_),
  .A2(_080_),
  .A3(_028_),
  .ZN(_081_)
);

NAND2_X1 _161_ (
  .A1(_030_),
  .A2(\coef[23] ),
  .ZN(_082_)
);

NAND2_X1 _162_ (
  .A1(_081_),
  .A2(_082_),
  .ZN(_003_)
);

NAND3_X1 _163_ (
  .A1(_056_),
  .A2(_058_),
  .A3(_038_),
  .ZN(_083_)
);

NAND3_X1 _164_ (
  .A1(_033_),
  .A2(_036_),
  .A3(_034_),
  .ZN(_084_)
);

NAND3_X1 _165_ (
  .A1(_065_),
  .A2(_048_),
  .A3(_084_),
  .ZN(_085_)
);

NAND3_X1 _166_ (
  .A1(_083_),
  .A2(_085_),
  .A3(_028_),
  .ZN(_086_)
);

NAND2_X1 _167_ (
  .A1(_030_),
  .A2(\coef[24] ),
  .ZN(_087_)
);

NAND2_X1 _168_ (
  .A1(_086_),
  .A2(_087_),
  .ZN(_004_)
);

NAND3_X1 _169_ (
  .A1(_078_),
  .A2(_069_),
  .A3(_048_),
  .ZN(_088_)
);

NAND3_X1 _170_ (
  .A1(_064_),
  .A2(_075_),
  .A3(_058_),
  .ZN(_089_)
);

NAND3_X1 _171_ (
  .A1(_088_),
  .A2(_089_),
  .A3(_028_),
  .ZN(_090_)
);

NAND2_X1 _172_ (
  .A1(_030_),
  .A2(\coef[25] ),
  .ZN(_091_)
);

NAND2_X1 _173_ (
  .A1(_090_),
  .A2(_091_),
  .ZN(_005_)
);

NAND3_X1 _174_ (
  .A1(_055_),
  .A2(_051_),
  .A3(_037_),
  .ZN(_092_)
);

NAND2_X1 _175_ (
  .A1(_056_),
  .A2(_092_),
  .ZN(_010_)
);

NAND2_X1 _176_ (
  .A1(_010_),
  .A2(_048_),
  .ZN(_011_)
);

NAND2_X1 _177_ (
  .A1(_062_),
  .A2(_047_),
  .ZN(_012_)
);

NAND2_X1 _178_ (
  .A1(_012_),
  .A2(_036_),
  .ZN(_013_)
);

NAND2_X1 _179_ (
  .A1(_035_),
  .A2(_046_),
  .ZN(_014_)
);

NAND3_X1 _180_ (
  .A1(_014_),
  .A2(_052_),
  .A3(_037_),
  .ZN(_015_)
);

NAND3_X1 _181_ (
  .A1(_013_),
  .A2(_015_),
  .A3(_058_),
  .ZN(_016_)
);

NAND3_X1 _182_ (
  .A1(_011_),
  .A2(_016_),
  .A3(_028_),
  .ZN(_017_)
);

NAND2_X1 _183_ (
  .A1(_030_),
  .A2(\coef[26] ),
  .ZN(_018_)
);

NAND2_X1 _184_ (
  .A1(_017_),
  .A2(_018_),
  .ZN(_006_)
);

NAND2_X1 _185_ (
  .A1(_030_),
  .A2(\coef[27] ),
  .ZN(_019_)
);

OAI21_X1 _186_ (
  .A(_028_),
  .B1(_043_),
  .B2(_048_),
  .ZN(_020_)
);

NAND3_X1 _187_ (
  .A1(_060_),
  .A2(_061_),
  .A3(_037_),
  .ZN(_021_)
);

AND3_X1 _188_ (
  .A1(_021_),
  .A2(_084_),
  .A3(_048_),
  .ZN(_022_)
);

OAI21_X1 _189_ (
  .A(_019_),
  .B1(_020_),
  .B2(_022_),
  .ZN(_007_)
);

NAND3_X1 _190_ (
  .A1(_064_),
  .A2(_079_),
  .A3(_048_),
  .ZN(_023_)
);

NAND3_X1 _191_ (
  .A1(_069_),
  .A2(_076_),
  .A3(_058_),
  .ZN(_024_)
);

NAND3_X1 _192_ (
  .A1(_023_),
  .A2(_024_),
  .A3(_028_),
  .ZN(_025_)
);

NAND2_X1 _193_ (
  .A1(_030_),
  .A2(\coef[28] ),
  .ZN(_026_)
);

NAND2_X1 _194_ (
  .A1(_025_),
  .A2(_026_),
  .ZN(_008_)
);

MUX2_X1 _195_ (
  .A(\coef[30] ),
  .B(_063_),
  .S(_027_),
  .Z(_009_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_101_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_100_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_099_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_098_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_097_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_096_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_095_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_094_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_102_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_093_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$32a02d514417e24bb09b7885b9c053483ac7784d\dctu

module \$paramod$37cd075c9fa8b3a4872c05f999800e89bc604dc4\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _196_ (
  .A(x[0]),
  .ZN(_178_)
);

INV_X1 _197_ (
  .A(x[1]),
  .ZN(_179_)
);

CLKBUF_X3 _198_ (
  .A(ena),
  .Z(_109_)
);

INV_X1 _199_ (
  .A(_109_),
  .ZN(_110_)
);

BUF_X8 _200_ (
  .A(x[2]),
  .Z(_111_)
);

INV_X8 _201_ (
  .A(_111_),
  .ZN(_112_)
);

NAND2_X4 _202_ (
  .A1(_112_),
  .A2(_180_),
  .ZN(_113_)
);

INV_X1 _203_ (
  .A(_194_),
  .ZN(_114_)
);

BUF_X32 _204_ (
  .A(_111_),
  .Z(_115_)
);

NAND2_X4 _205_ (
  .A1(_114_),
  .A2(_115_),
  .ZN(_116_)
);

BUF_X8 _206_ (
  .A(y[0]),
  .Z(_117_)
);

BUF_X16 _207_ (
  .A(_117_),
  .Z(_118_)
);

NAND3_X4 _208_ (
  .A1(_113_),
  .A2(_116_),
  .A3(_118_),
  .ZN(_119_)
);

INV_X1 _209_ (
  .A(_181_),
  .ZN(_120_)
);

NAND2_X4 _210_ (
  .A1(_112_),
  .A2(_120_),
  .ZN(_121_)
);

NAND2_X2 _211_ (
  .A1(_111_),
  .A2(_181_),
  .ZN(_122_)
);

NAND2_X4 _212_ (
  .A1(_121_),
  .A2(_122_),
  .ZN(_123_)
);

OAI21_X2 _213_ (
  .A(_119_),
  .B1(_118_),
  .B2(_123_),
  .ZN(_124_)
);

BUF_X4 _214_ (
  .A(y[1]),
  .Z(_125_)
);

INV_X2 _215_ (
  .A(_125_),
  .ZN(_126_)
);

BUF_X4 _216_ (
  .A(_126_),
  .Z(_127_)
);

NAND2_X1 _217_ (
  .A1(_124_),
  .A2(_127_),
  .ZN(_128_)
);

NAND2_X2 _218_ (
  .A1(_117_),
  .A2(x[1]),
  .ZN(_129_)
);

NAND2_X1 _219_ (
  .A1(_129_),
  .A2(_125_),
  .ZN(_130_)
);

NAND2_X4 _220_ (
  .A1(_112_),
  .A2(_188_),
  .ZN(_131_)
);

INV_X1 _221_ (
  .A(_186_),
  .ZN(_132_)
);

NAND2_X4 _222_ (
  .A1(_132_),
  .A2(_115_),
  .ZN(_133_)
);

NAND2_X2 _223_ (
  .A1(_131_),
  .A2(_133_),
  .ZN(_134_)
);

INV_X16 _224_ (
  .A(_117_),
  .ZN(_135_)
);

BUF_X16 _225_ (
  .A(_135_),
  .Z(_136_)
);

AOI21_X2 _226_ (
  .A(_130_),
  .B1(_134_),
  .B2(_136_),
  .ZN(_137_)
);

BUF_X2 _227_ (
  .A(y[2]),
  .Z(_138_)
);

INV_X1 _228_ (
  .A(_138_),
  .ZN(_139_)
);

BUF_X4 _229_ (
  .A(_139_),
  .Z(_140_)
);

NOR2_X2 _230_ (
  .A1(_137_),
  .A2(_140_),
  .ZN(_141_)
);

AOI21_X2 _231_ (
  .A(_110_),
  .B1(_128_),
  .B2(_141_),
  .ZN(_142_)
);

INV_X1 _232_ (
  .A(_182_),
  .ZN(_143_)
);

NAND2_X2 _233_ (
  .A1(_112_),
  .A2(_143_),
  .ZN(_144_)
);

NAND2_X4 _234_ (
  .A1(_115_),
  .A2(_192_),
  .ZN(_145_)
);

NAND3_X2 _235_ (
  .A1(_144_),
  .A2(_136_),
  .A3(_145_),
  .ZN(_146_)
);

INV_X1 _236_ (
  .A(_123_),
  .ZN(_147_)
);

OAI21_X1 _237_ (
  .A(_146_),
  .B1(_147_),
  .B2(_136_),
  .ZN(_148_)
);

BUF_X2 _238_ (
  .A(_125_),
  .Z(_149_)
);

NAND2_X1 _239_ (
  .A1(_148_),
  .A2(_149_),
  .ZN(_150_)
);

INV_X1 _240_ (
  .A(_190_),
  .ZN(_151_)
);

NAND2_X4 _241_ (
  .A1(_112_),
  .A2(_151_),
  .ZN(_152_)
);

NAND2_X4 _242_ (
  .A1(_115_),
  .A2(_184_),
  .ZN(_153_)
);

NAND2_X2 _243_ (
  .A1(_152_),
  .A2(_153_),
  .ZN(_154_)
);

NAND2_X1 _244_ (
  .A1(_154_),
  .A2(_118_),
  .ZN(_155_)
);

NAND2_X1 _245_ (
  .A1(_135_),
  .A2(_179_),
  .ZN(_156_)
);

NAND3_X1 _246_ (
  .A1(_155_),
  .A2(_127_),
  .A3(_156_),
  .ZN(_157_)
);

NAND3_X1 _247_ (
  .A1(_150_),
  .A2(_140_),
  .A3(_157_),
  .ZN(_158_)
);

NAND2_X1 _248_ (
  .A1(_142_),
  .A2(_158_),
  .ZN(_159_)
);

NAND2_X1 _249_ (
  .A1(_110_),
  .A2(\coef[21] ),
  .ZN(_160_)
);

NAND2_X1 _250_ (
  .A1(_159_),
  .A2(_160_),
  .ZN(_000_)
);

NAND3_X1 _251_ (
  .A1(_131_),
  .A2(_133_),
  .A3(_136_),
  .ZN(_161_)
);

NAND3_X2 _252_ (
  .A1(_144_),
  .A2(_118_),
  .A3(_145_),
  .ZN(_162_)
);

NAND3_X1 _253_ (
  .A1(_161_),
  .A2(_162_),
  .A3(_126_),
  .ZN(_163_)
);

NAND3_X1 _254_ (
  .A1(_156_),
  .A2(_149_),
  .A3(_129_),
  .ZN(_164_)
);

NAND3_X1 _255_ (
  .A1(_163_),
  .A2(_138_),
  .A3(_164_),
  .ZN(_165_)
);

NAND3_X2 _256_ (
  .A1(_113_),
  .A2(_116_),
  .A3(_136_),
  .ZN(_166_)
);

NAND3_X1 _257_ (
  .A1(_152_),
  .A2(_118_),
  .A3(_153_),
  .ZN(_167_)
);

NAND3_X1 _258_ (
  .A1(_166_),
  .A2(_167_),
  .A3(_149_),
  .ZN(_168_)
);

NAND3_X1 _259_ (
  .A1(_156_),
  .A2(_126_),
  .A3(_129_),
  .ZN(_009_)
);

NAND3_X1 _260_ (
  .A1(_168_),
  .A2(_140_),
  .A3(_009_),
  .ZN(_010_)
);

NAND2_X1 _261_ (
  .A1(_165_),
  .A2(_010_),
  .ZN(_011_)
);

NAND2_X1 _262_ (
  .A1(_011_),
  .A2(_109_),
  .ZN(_012_)
);

NAND2_X1 _263_ (
  .A1(_110_),
  .A2(\coef[23] ),
  .ZN(_013_)
);

NAND2_X1 _264_ (
  .A1(_012_),
  .A2(_013_),
  .ZN(_001_)
);

NAND2_X2 _265_ (
  .A1(_112_),
  .A2(_186_),
  .ZN(_014_)
);

INV_X1 _266_ (
  .A(_188_),
  .ZN(_015_)
);

NAND2_X4 _267_ (
  .A1(_015_),
  .A2(_115_),
  .ZN(_016_)
);

NAND2_X2 _268_ (
  .A1(_014_),
  .A2(_016_),
  .ZN(_017_)
);

NAND2_X4 _269_ (
  .A1(_017_),
  .A2(_118_),
  .ZN(_018_)
);

NOR2_X2 _270_ (
  .A1(_115_),
  .A2(_117_),
  .ZN(_019_)
);

INV_X1 _271_ (
  .A(_019_),
  .ZN(_020_)
);

NAND3_X1 _272_ (
  .A1(_018_),
  .A2(_149_),
  .A3(_020_),
  .ZN(_021_)
);

NAND3_X4 _273_ (
  .A1(_131_),
  .A2(_133_),
  .A3(_117_),
  .ZN(_022_)
);

NAND3_X1 _274_ (
  .A1(_022_),
  .A2(_126_),
  .A3(_156_),
  .ZN(_023_)
);

NAND3_X1 _275_ (
  .A1(_021_),
  .A2(_023_),
  .A3(_140_),
  .ZN(_024_)
);

INV_X1 _276_ (
  .A(_184_),
  .ZN(_025_)
);

NAND2_X1 _277_ (
  .A1(_112_),
  .A2(_025_),
  .ZN(_026_)
);

NAND2_X4 _278_ (
  .A1(_115_),
  .A2(_190_),
  .ZN(_027_)
);

NAND2_X2 _279_ (
  .A1(_026_),
  .A2(_027_),
  .ZN(_028_)
);

NAND2_X2 _280_ (
  .A1(_028_),
  .A2(_136_),
  .ZN(_029_)
);

NAND2_X4 _281_ (
  .A1(_115_),
  .A2(_117_),
  .ZN(_030_)
);

NAND3_X1 _282_ (
  .A1(_029_),
  .A2(_126_),
  .A3(_030_),
  .ZN(_031_)
);

NAND3_X4 _283_ (
  .A1(_152_),
  .A2(_135_),
  .A3(_153_),
  .ZN(_032_)
);

NAND3_X1 _284_ (
  .A1(_032_),
  .A2(_125_),
  .A3(_129_),
  .ZN(_033_)
);

NAND3_X1 _285_ (
  .A1(_031_),
  .A2(_033_),
  .A3(_138_),
  .ZN(_034_)
);

NAND2_X1 _286_ (
  .A1(_024_),
  .A2(_034_),
  .ZN(_035_)
);

NAND2_X1 _287_ (
  .A1(_035_),
  .A2(_109_),
  .ZN(_036_)
);

NAND2_X1 _288_ (
  .A1(_110_),
  .A2(\coef[24] ),
  .ZN(_037_)
);

NAND2_X2 _289_ (
  .A1(_036_),
  .A2(_037_),
  .ZN(_002_)
);

OAI21_X1 _290_ (
  .A(_125_),
  .B1(_135_),
  .B2(x[0]),
  .ZN(_038_)
);

INV_X1 _291_ (
  .A(_038_),
  .ZN(_039_)
);

AOI21_X1 _292_ (
  .A(_138_),
  .B1(_039_),
  .B2(_156_),
  .ZN(_040_)
);

INV_X1 _293_ (
  .A(_030_),
  .ZN(_041_)
);

AOI21_X1 _294_ (
  .A(_041_),
  .B1(_147_),
  .B2(_136_),
  .ZN(_042_)
);

OAI21_X1 _295_ (
  .A(_040_),
  .B1(_042_),
  .B2(_149_),
  .ZN(_043_)
);

NAND2_X1 _296_ (
  .A1(_129_),
  .A2(_126_),
  .ZN(_044_)
);

INV_X1 _297_ (
  .A(_044_),
  .ZN(_045_)
);

NOR2_X1 _298_ (
  .A1(_178_),
  .A2(_117_),
  .ZN(_046_)
);

INV_X1 _299_ (
  .A(_046_),
  .ZN(_047_)
);

AOI21_X1 _300_ (
  .A(_139_),
  .B1(_045_),
  .B2(_047_),
  .ZN(_048_)
);

AOI21_X1 _301_ (
  .A(_019_),
  .B1(_123_),
  .B2(_118_),
  .ZN(_049_)
);

OAI21_X1 _302_ (
  .A(_048_),
  .B1(_049_),
  .B2(_127_),
  .ZN(_050_)
);

NAND3_X1 _303_ (
  .A1(_043_),
  .A2(_050_),
  .A3(_109_),
  .ZN(_051_)
);

NAND2_X1 _304_ (
  .A1(_110_),
  .A2(\coef[10] ),
  .ZN(_052_)
);

NAND2_X1 _305_ (
  .A1(_051_),
  .A2(_052_),
  .ZN(_003_)
);

NOR2_X1 _306_ (
  .A1(_109_),
  .A2(\coef[26] ),
  .ZN(_053_)
);

AOI21_X1 _307_ (
  .A(_140_),
  .B1(_166_),
  .B2(_045_),
  .ZN(_054_)
);

NAND3_X1 _308_ (
  .A1(_121_),
  .A2(_118_),
  .A3(_122_),
  .ZN(_055_)
);

NAND3_X1 _309_ (
  .A1(_146_),
  .A2(_055_),
  .A3(_149_),
  .ZN(_056_)
);

AOI21_X1 _310_ (
  .A(_110_),
  .B1(_054_),
  .B2(_056_),
  .ZN(_057_)
);

NAND2_X2 _311_ (
  .A1(_123_),
  .A2(_136_),
  .ZN(_058_)
);

NAND2_X1 _312_ (
  .A1(_058_),
  .A2(_119_),
  .ZN(_059_)
);

NAND2_X1 _313_ (
  .A1(_059_),
  .A2(_127_),
  .ZN(_060_)
);

NAND2_X1 _314_ (
  .A1(_162_),
  .A2(_156_),
  .ZN(_061_)
);

NAND2_X1 _315_ (
  .A1(_061_),
  .A2(_149_),
  .ZN(_062_)
);

NAND2_X1 _316_ (
  .A1(_060_),
  .A2(_062_),
  .ZN(_063_)
);

NAND2_X1 _317_ (
  .A1(_063_),
  .A2(_140_),
  .ZN(_064_)
);

AOI21_X2 _318_ (
  .A(_053_),
  .B1(_057_),
  .B2(_064_),
  .ZN(_004_)
);

NAND2_X1 _319_ (
  .A1(_112_),
  .A2(_192_),
  .ZN(_065_)
);

NAND2_X2 _320_ (
  .A1(_143_),
  .A2(_115_),
  .ZN(_066_)
);

NAND3_X2 _321_ (
  .A1(_065_),
  .A2(_066_),
  .A3(_118_),
  .ZN(_067_)
);

NAND3_X1 _322_ (
  .A1(_067_),
  .A2(_127_),
  .A3(_020_),
  .ZN(_068_)
);

NAND2_X1 _323_ (
  .A1(_029_),
  .A2(_039_),
  .ZN(_069_)
);

NAND3_X1 _324_ (
  .A1(_068_),
  .A2(_140_),
  .A3(_069_),
  .ZN(_070_)
);

NAND2_X1 _325_ (
  .A1(_112_),
  .A2(_114_),
  .ZN(_071_)
);

NAND2_X4 _326_ (
  .A1(_115_),
  .A2(_180_),
  .ZN(_072_)
);

NAND3_X2 _327_ (
  .A1(_071_),
  .A2(_136_),
  .A3(_072_),
  .ZN(_073_)
);

NAND2_X4 _328_ (
  .A1(_030_),
  .A2(_125_),
  .ZN(_074_)
);

INV_X2 _329_ (
  .A(_074_),
  .ZN(_075_)
);

AOI21_X2 _330_ (
  .A(_139_),
  .B1(_073_),
  .B2(_075_),
  .ZN(_076_)
);

NAND3_X1 _331_ (
  .A1(_018_),
  .A2(_126_),
  .A3(_047_),
  .ZN(_077_)
);

NAND2_X1 _332_ (
  .A1(_076_),
  .A2(_077_),
  .ZN(_078_)
);

NAND3_X1 _333_ (
  .A1(_070_),
  .A2(_109_),
  .A3(_078_),
  .ZN(_079_)
);

OR2_X1 _334_ (
  .A1(\coef[13] ),
  .A2(_109_),
  .ZN(_080_)
);

AND2_X2 _335_ (
  .A1(_079_),
  .A2(_080_),
  .ZN(_005_)
);

NAND3_X1 _336_ (
  .A1(_071_),
  .A2(_118_),
  .A3(_072_),
  .ZN(_081_)
);

NAND3_X1 _337_ (
  .A1(_029_),
  .A2(_081_),
  .A3(_126_),
  .ZN(_082_)
);

NAND3_X1 _338_ (
  .A1(_119_),
  .A2(_032_),
  .A3(_125_),
  .ZN(_083_)
);

NAND3_X1 _339_ (
  .A1(_082_),
  .A2(_083_),
  .A3(_138_),
  .ZN(_084_)
);

NAND3_X1 _340_ (
  .A1(_065_),
  .A2(_066_),
  .A3(_136_),
  .ZN(_085_)
);

NAND3_X2 _341_ (
  .A1(_018_),
  .A2(_085_),
  .A3(_149_),
  .ZN(_086_)
);

NAND3_X1 _342_ (
  .A1(_022_),
  .A2(_146_),
  .A3(_126_),
  .ZN(_087_)
);

NAND3_X1 _343_ (
  .A1(_086_),
  .A2(_087_),
  .A3(_140_),
  .ZN(_088_)
);

NAND2_X1 _344_ (
  .A1(_084_),
  .A2(_088_),
  .ZN(_089_)
);

NAND2_X1 _345_ (
  .A1(_089_),
  .A2(_109_),
  .ZN(_090_)
);

NAND2_X1 _346_ (
  .A1(_110_),
  .A2(\coef[28] ),
  .ZN(_091_)
);

NAND2_X1 _347_ (
  .A1(_090_),
  .A2(_091_),
  .ZN(_006_)
);

NAND2_X1 _348_ (
  .A1(_022_),
  .A2(_073_),
  .ZN(_092_)
);

NAND2_X1 _349_ (
  .A1(_092_),
  .A2(_127_),
  .ZN(_093_)
);

NAND2_X1 _350_ (
  .A1(_058_),
  .A2(_075_),
  .ZN(_094_)
);

NAND3_X1 _351_ (
  .A1(_093_),
  .A2(_140_),
  .A3(_094_),
  .ZN(_095_)
);

NAND2_X1 _352_ (
  .A1(_067_),
  .A2(_032_),
  .ZN(_096_)
);

NAND2_X1 _353_ (
  .A1(_096_),
  .A2(_149_),
  .ZN(_097_)
);

NAND3_X1 _354_ (
  .A1(_055_),
  .A2(_127_),
  .A3(_020_),
  .ZN(_098_)
);

NAND3_X1 _355_ (
  .A1(_097_),
  .A2(_098_),
  .A3(_138_),
  .ZN(_099_)
);

NAND3_X1 _356_ (
  .A1(_095_),
  .A2(_099_),
  .A3(_109_),
  .ZN(_100_)
);

NAND2_X1 _357_ (
  .A1(_110_),
  .A2(\coef[29] ),
  .ZN(_101_)
);

NAND2_X1 _358_ (
  .A1(_100_),
  .A2(_101_),
  .ZN(_007_)
);

NOR2_X1 _359_ (
  .A1(_109_),
  .A2(\coef[30] ),
  .ZN(_102_)
);

NAND3_X1 _360_ (
  .A1(_022_),
  .A2(_032_),
  .A3(_127_),
  .ZN(_103_)
);

AOI21_X1 _361_ (
  .A(_138_),
  .B1(_134_),
  .B2(_149_),
  .ZN(_104_)
);

AOI21_X1 _362_ (
  .A(_110_),
  .B1(_103_),
  .B2(_104_),
  .ZN(_105_)
);

AOI21_X1 _363_ (
  .A(_140_),
  .B1(_154_),
  .B2(_127_),
  .ZN(_106_)
);

NAND2_X1 _364_ (
  .A1(_022_),
  .A2(_032_),
  .ZN(_107_)
);

OAI21_X1 _365_ (
  .A(_106_),
  .B1(_107_),
  .B2(_127_),
  .ZN(_108_)
);

AOI21_X1 _366_ (
  .A(_102_),
  .B1(_105_),
  .B2(_108_),
  .ZN(_008_)
);

HA_X1 _367_ (
  .A(_178_),
  .B(_179_),
  .CO(_180_),
  .S(_181_)
);

HA_X1 _368_ (
  .A(_178_),
  .B(_179_),
  .CO(_182_),
  .S(_183_)
);

HA_X1 _369_ (
  .A(_178_),
  .B(x[1]),
  .CO(_184_),
  .S(_185_)
);

HA_X1 _370_ (
  .A(_178_),
  .B(x[1]),
  .CO(_186_),
  .S(_187_)
);

HA_X1 _371_ (
  .A(x[0]),
  .B(_179_),
  .CO(_188_),
  .S(_189_)
);

HA_X1 _372_ (
  .A(x[0]),
  .B(_179_),
  .CO(_190_),
  .S(_191_)
);

HA_X1 _373_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_192_),
  .S(_193_)
);

HA_X1 _374_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_194_),
  .S(_195_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_177_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_176_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_175_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_174_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_173_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_172_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_171_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_170_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_169_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$37cd075c9fa8b3a4872c05f999800e89bc604dc4\dctu

module \$paramod$3b47752d19f391915a818678f43c9a51f524cc48\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _11_ (
  .A(y[1]),
  .ZN(_04_)
);

INV_X1 _12_ (
  .A(y[0]),
  .ZN(_05_)
);

NAND2_X1 _13_ (
  .A1(_04_),
  .A2(_05_),
  .ZN(_06_)
);

NAND2_X1 _14_ (
  .A1(y[1]),
  .A2(y[0]),
  .ZN(_07_)
);

NAND3_X1 _15_ (
  .A1(_06_),
  .A2(ena),
  .A3(_07_),
  .ZN(_01_)
);

INV_X1 _16_ (
  .A(ena),
  .ZN(_02_)
);

NAND2_X1 _17_ (
  .A1(_02_),
  .A2(\coef[30] ),
  .ZN(_03_)
);

NAND2_X1 _18_ (
  .A1(_01_),
  .A2(_03_),
  .ZN(_00_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_08_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_47974  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , _09_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_}),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$3b47752d19f391915a818678f43c9a51f524cc48\dctu

module \$paramod$44a044575968c599376fc32b4d9ee49faea5711d\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _090_ (
  .A(x[0]),
  .ZN(_072_)
);

INV_X1 _091_ (
  .A(x[1]),
  .ZN(_073_)
);

BUF_X8 _092_ (
  .A(x[2]),
  .Z(_008_)
);

NOR2_X1 _093_ (
  .A1(_008_),
  .A2(_078_),
  .ZN(_009_)
);

AOI21_X1 _094_ (
  .A(_009_),
  .B1(_084_),
  .B2(_008_),
  .ZN(_010_)
);

INV_X2 _095_ (
  .A(y[0]),
  .ZN(_011_)
);

INV_X1 _096_ (
  .A(y[1]),
  .ZN(_012_)
);

NAND2_X2 _097_ (
  .A1(_011_),
  .A2(_012_),
  .ZN(_013_)
);

NAND2_X1 _098_ (
  .A1(y[0]),
  .A2(y[1]),
  .ZN(_014_)
);

NAND2_X4 _099_ (
  .A1(_013_),
  .A2(_014_),
  .ZN(_015_)
);

INV_X2 _100_ (
  .A(_015_),
  .ZN(_016_)
);

NAND2_X1 _101_ (
  .A1(_010_),
  .A2(_016_),
  .ZN(_017_)
);

BUF_X1 _102_ (
  .A(ena),
  .Z(_018_)
);

BUF_X4 _103_ (
  .A(_018_),
  .Z(_019_)
);

INV_X8 _104_ (
  .A(_008_),
  .ZN(_020_)
);

OR2_X4 _105_ (
  .A1(_020_),
  .A2(_082_),
  .ZN(_021_)
);

NAND2_X1 _106_ (
  .A1(_020_),
  .A2(_080_),
  .ZN(_022_)
);

NAND3_X1 _107_ (
  .A1(_015_),
  .A2(_021_),
  .A3(_022_),
  .ZN(_023_)
);

NAND3_X1 _108_ (
  .A1(_017_),
  .A2(_019_),
  .A3(_023_),
  .ZN(_024_)
);

INV_X1 _109_ (
  .A(_018_),
  .ZN(_025_)
);

NAND2_X1 _110_ (
  .A1(_025_),
  .A2(\coef[21] ),
  .ZN(_026_)
);

NAND2_X1 _111_ (
  .A1(_024_),
  .A2(_026_),
  .ZN(_000_)
);

XNOR2_X2 _112_ (
  .A(_015_),
  .B(_073_),
  .ZN(_027_)
);

NAND2_X2 _113_ (
  .A1(_027_),
  .A2(_019_),
  .ZN(_028_)
);

INV_X1 _114_ (
  .A(\coef[22] ),
  .ZN(_029_)
);

OAI21_X2 _115_ (
  .A(_028_),
  .B1(_019_),
  .B2(_029_),
  .ZN(_001_)
);

NAND2_X1 _116_ (
  .A1(_015_),
  .A2(_008_),
  .ZN(_030_)
);

NAND3_X1 _117_ (
  .A1(_013_),
  .A2(_020_),
  .A3(_014_),
  .ZN(_031_)
);

NAND3_X1 _118_ (
  .A1(_030_),
  .A2(_031_),
  .A3(_019_),
  .ZN(_032_)
);

INV_X1 _119_ (
  .A(\coef[23] ),
  .ZN(_033_)
);

OAI21_X1 _120_ (
  .A(_032_),
  .B1(_019_),
  .B2(_033_),
  .ZN(_002_)
);

NOR2_X1 _121_ (
  .A1(_018_),
  .A2(\coef[14] ),
  .ZN(_034_)
);

AOI21_X2 _122_ (
  .A(_034_),
  .B1(_027_),
  .B2(_019_),
  .ZN(_003_)
);

NAND2_X1 _123_ (
  .A1(_008_),
  .A2(_088_),
  .ZN(_035_)
);

INV_X1 _124_ (
  .A(_074_),
  .ZN(_036_)
);

NAND2_X1 _125_ (
  .A1(_020_),
  .A2(_036_),
  .ZN(_037_)
);

NAND3_X1 _126_ (
  .A1(_016_),
  .A2(_035_),
  .A3(_037_),
  .ZN(_038_)
);

OR2_X4 _127_ (
  .A1(_020_),
  .A2(_086_),
  .ZN(_039_)
);

NAND2_X1 _128_ (
  .A1(_020_),
  .A2(_076_),
  .ZN(_040_)
);

NAND3_X1 _129_ (
  .A1(_015_),
  .A2(_039_),
  .A3(_040_),
  .ZN(_041_)
);

NAND3_X1 _130_ (
  .A1(_038_),
  .A2(_019_),
  .A3(_041_),
  .ZN(_042_)
);

NAND2_X1 _131_ (
  .A1(_025_),
  .A2(\coef[13] ),
  .ZN(_043_)
);

NAND2_X1 _132_ (
  .A1(_042_),
  .A2(_043_),
  .ZN(_004_)
);

NOR2_X1 _133_ (
  .A1(_008_),
  .A2(_086_),
  .ZN(_044_)
);

AOI21_X1 _134_ (
  .A(_044_),
  .B1(_076_),
  .B2(_008_),
  .ZN(_045_)
);

NAND2_X1 _135_ (
  .A1(_045_),
  .A2(_016_),
  .ZN(_046_)
);

NAND2_X1 _136_ (
  .A1(_036_),
  .A2(_008_),
  .ZN(_047_)
);

NAND2_X1 _137_ (
  .A1(_020_),
  .A2(_088_),
  .ZN(_048_)
);

NAND3_X1 _138_ (
  .A1(_015_),
  .A2(_047_),
  .A3(_048_),
  .ZN(_049_)
);

NAND3_X1 _139_ (
  .A1(_046_),
  .A2(_019_),
  .A3(_049_),
  .ZN(_050_)
);

NAND2_X1 _140_ (
  .A1(_025_),
  .A2(\coef[28] ),
  .ZN(_051_)
);

NAND2_X1 _141_ (
  .A1(_050_),
  .A2(_051_),
  .ZN(_005_)
);

INV_X1 _142_ (
  .A(_075_),
  .ZN(_052_)
);

NAND3_X1 _143_ (
  .A1(_030_),
  .A2(_031_),
  .A3(_052_),
  .ZN(_053_)
);

NAND2_X4 _144_ (
  .A1(_020_),
  .A2(_011_),
  .ZN(_054_)
);

NAND2_X1 _145_ (
  .A1(_008_),
  .A2(y[0]),
  .ZN(_055_)
);

NAND2_X1 _146_ (
  .A1(_054_),
  .A2(_055_),
  .ZN(_056_)
);

NAND2_X1 _147_ (
  .A1(_056_),
  .A2(_012_),
  .ZN(_057_)
);

NAND3_X1 _148_ (
  .A1(_054_),
  .A2(y[1]),
  .A3(_055_),
  .ZN(_058_)
);

NAND3_X1 _149_ (
  .A1(_057_),
  .A2(_058_),
  .A3(_075_),
  .ZN(_059_)
);

NAND3_X1 _150_ (
  .A1(_053_),
  .A2(_059_),
  .A3(_019_),
  .ZN(_060_)
);

NAND2_X1 _151_ (
  .A1(_025_),
  .A2(\coef[15] ),
  .ZN(_061_)
);

NAND2_X1 _152_ (
  .A1(_060_),
  .A2(_061_),
  .ZN(_006_)
);

NOR2_X1 _153_ (
  .A1(_018_),
  .A2(\coef[12] ),
  .ZN(_062_)
);

XNOR2_X1 _154_ (
  .A(_015_),
  .B(_072_),
  .ZN(_063_)
);

AOI21_X2 _155_ (
  .A(_062_),
  .B1(_063_),
  .B2(_019_),
  .ZN(_007_)
);

HA_X1 _156_ (
  .A(_072_),
  .B(_073_),
  .CO(_074_),
  .S(_075_)
);

HA_X1 _157_ (
  .A(_072_),
  .B(_073_),
  .CO(_076_),
  .S(_077_)
);

HA_X1 _158_ (
  .A(_072_),
  .B(x[1]),
  .CO(_078_),
  .S(_079_)
);

HA_X1 _159_ (
  .A(_072_),
  .B(x[1]),
  .CO(_080_),
  .S(_081_)
);

HA_X1 _160_ (
  .A(x[0]),
  .B(_073_),
  .CO(_082_),
  .S(_083_)
);

HA_X1 _161_ (
  .A(x[0]),
  .B(_073_),
  .CO(_084_),
  .S(_085_)
);

HA_X1 _162_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_086_),
  .S(_087_)
);

HA_X1 _163_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_088_),
  .S(_089_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_071_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_070_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_069_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_068_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_067_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_066_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_065_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_064_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$44a044575968c599376fc32b4d9ee49faea5711d\dctu

module \$paramod$29130e85acc43116076719ea36da8d59b7490cc4\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _183_ (
  .A(x[1]),
  .ZN(_166_)
);

INV_X1 _184_ (
  .A(x[0]),
  .ZN(_165_)
);

CLKBUF_X2 _185_ (
  .A(y[2]),
  .Z(_097_)
);

BUF_X4 _186_ (
  .A(x[2]),
  .Z(_098_)
);

INV_X4 _187_ (
  .A(_098_),
  .ZN(_099_)
);

NAND2_X4 _188_ (
  .A1(_099_),
  .A2(_171_),
  .ZN(_100_)
);

INV_X1 _189_ (
  .A(_177_),
  .ZN(_101_)
);

BUF_X16 _190_ (
  .A(_098_),
  .Z(_102_)
);

NAND2_X4 _191_ (
  .A1(_101_),
  .A2(_102_),
  .ZN(_103_)
);

NAND2_X4 _192_ (
  .A1(_100_),
  .A2(_103_),
  .ZN(_104_)
);

BUF_X8 _193_ (
  .A(y[0]),
  .Z(_105_)
);

INV_X8 _194_ (
  .A(_105_),
  .ZN(_106_)
);

BUF_X8 _195_ (
  .A(_106_),
  .Z(_107_)
);

NAND2_X2 _196_ (
  .A1(_104_),
  .A2(_107_),
  .ZN(_108_)
);

BUF_X4 _197_ (
  .A(y[1]),
  .Z(_109_)
);

OAI21_X2 _198_ (
  .A(_109_),
  .B1(_106_),
  .B2(_165_),
  .ZN(_110_)
);

INV_X1 _199_ (
  .A(_110_),
  .ZN(_111_)
);

AOI21_X2 _200_ (
  .A(_097_),
  .B1(_108_),
  .B2(_111_),
  .ZN(_112_)
);

BUF_X2 _201_ (
  .A(_109_),
  .Z(_113_)
);

NAND2_X2 _202_ (
  .A1(_099_),
  .A2(_179_),
  .ZN(_114_)
);

INV_X1 _203_ (
  .A(_169_),
  .ZN(_115_)
);

NAND2_X4 _204_ (
  .A1(_115_),
  .A2(_102_),
  .ZN(_116_)
);

BUF_X8 _205_ (
  .A(_105_),
  .Z(_117_)
);

NAND3_X2 _206_ (
  .A1(_114_),
  .A2(_116_),
  .A3(_117_),
  .ZN(_118_)
);

NOR2_X4 _207_ (
  .A1(_102_),
  .A2(_105_),
  .ZN(_119_)
);

INV_X1 _208_ (
  .A(_119_),
  .ZN(_120_)
);

AND2_X2 _209_ (
  .A1(_118_),
  .A2(_120_),
  .ZN(_121_)
);

OAI21_X2 _210_ (
  .A(_112_),
  .B1(_113_),
  .B2(_121_),
  .ZN(_122_)
);

INV_X1 _211_ (
  .A(_181_),
  .ZN(_123_)
);

NAND2_X2 _212_ (
  .A1(_099_),
  .A2(_123_),
  .ZN(_124_)
);

NAND2_X4 _213_ (
  .A1(_102_),
  .A2(_167_),
  .ZN(_125_)
);

NAND3_X1 _214_ (
  .A1(_124_),
  .A2(_106_),
  .A3(_125_),
  .ZN(_126_)
);

INV_X1 _215_ (
  .A(_126_),
  .ZN(_127_)
);

NAND2_X4 _216_ (
  .A1(_102_),
  .A2(_105_),
  .ZN(_128_)
);

INV_X1 _217_ (
  .A(_128_),
  .ZN(_129_)
);

OAI21_X1 _218_ (
  .A(_113_),
  .B1(_127_),
  .B2(_129_),
  .ZN(_130_)
);

INV_X1 _219_ (
  .A(_097_),
  .ZN(_131_)
);

BUF_X4 _220_ (
  .A(_131_),
  .Z(_132_)
);

INV_X1 _221_ (
  .A(_173_),
  .ZN(_133_)
);

NAND2_X2 _222_ (
  .A1(_099_),
  .A2(_133_),
  .ZN(_134_)
);

NAND2_X4 _223_ (
  .A1(_102_),
  .A2(_175_),
  .ZN(_135_)
);

NAND2_X2 _224_ (
  .A1(_134_),
  .A2(_135_),
  .ZN(_136_)
);

NAND2_X1 _225_ (
  .A1(_136_),
  .A2(_117_),
  .ZN(_137_)
);

NOR2_X2 _226_ (
  .A1(_105_),
  .A2(x[0]),
  .ZN(_138_)
);

NOR2_X1 _227_ (
  .A1(_138_),
  .A2(_109_),
  .ZN(_139_)
);

AOI21_X1 _228_ (
  .A(_132_),
  .B1(_137_),
  .B2(_139_),
  .ZN(_140_)
);

NAND2_X1 _229_ (
  .A1(_130_),
  .A2(_140_),
  .ZN(_141_)
);

BUF_X2 _230_ (
  .A(ena),
  .Z(_142_)
);

NAND3_X1 _231_ (
  .A1(_122_),
  .A2(_141_),
  .A3(_142_),
  .ZN(_143_)
);

INV_X1 _232_ (
  .A(_142_),
  .ZN(_144_)
);

NAND2_X1 _233_ (
  .A1(_144_),
  .A2(\coef[21] ),
  .ZN(_145_)
);

NAND2_X1 _234_ (
  .A1(_143_),
  .A2(_145_),
  .ZN(_000_)
);

OAI21_X1 _235_ (
  .A(_110_),
  .B1(_113_),
  .B2(_129_),
  .ZN(_146_)
);

NAND3_X1 _236_ (
  .A1(_134_),
  .A2(_106_),
  .A3(_135_),
  .ZN(_147_)
);

NAND3_X1 _237_ (
  .A1(_146_),
  .A2(_132_),
  .A3(_147_),
  .ZN(_148_)
);

INV_X1 _238_ (
  .A(_109_),
  .ZN(_149_)
);

NOR2_X1 _239_ (
  .A1(_119_),
  .A2(_149_),
  .ZN(_150_)
);

OR2_X2 _240_ (
  .A1(_150_),
  .A2(_139_),
  .ZN(_151_)
);

NAND3_X4 _241_ (
  .A1(_100_),
  .A2(_103_),
  .A3(_105_),
  .ZN(_152_)
);

NAND3_X1 _242_ (
  .A1(_151_),
  .A2(_097_),
  .A3(_152_),
  .ZN(_153_)
);

NAND3_X1 _243_ (
  .A1(_148_),
  .A2(_153_),
  .A3(_142_),
  .ZN(_154_)
);

INV_X1 _244_ (
  .A(\coef[23] ),
  .ZN(_155_)
);

OAI21_X1 _245_ (
  .A(_154_),
  .B1(_142_),
  .B2(_155_),
  .ZN(_001_)
);

XNOR2_X2 _246_ (
  .A(_098_),
  .B(_168_),
  .ZN(_009_)
);

NAND2_X2 _247_ (
  .A1(_009_),
  .A2(_107_),
  .ZN(_010_)
);

NAND2_X1 _248_ (
  .A1(_128_),
  .A2(_109_),
  .ZN(_011_)
);

INV_X1 _249_ (
  .A(_011_),
  .ZN(_012_)
);

AOI21_X4 _250_ (
  .A(_131_),
  .B1(_010_),
  .B2(_012_),
  .ZN(_013_)
);

NAND2_X2 _251_ (
  .A1(_099_),
  .A2(_115_),
  .ZN(_014_)
);

NAND2_X4 _252_ (
  .A1(_102_),
  .A2(_179_),
  .ZN(_015_)
);

NAND3_X2 _253_ (
  .A1(_014_),
  .A2(_106_),
  .A3(_015_),
  .ZN(_016_)
);

NAND2_X1 _254_ (
  .A1(_152_),
  .A2(_016_),
  .ZN(_017_)
);

BUF_X4 _255_ (
  .A(_149_),
  .Z(_018_)
);

NAND2_X1 _256_ (
  .A1(_017_),
  .A2(_018_),
  .ZN(_019_)
);

AOI21_X2 _257_ (
  .A(_144_),
  .B1(_013_),
  .B2(_019_),
  .ZN(_020_)
);

NAND2_X2 _258_ (
  .A1(_099_),
  .A2(_167_),
  .ZN(_021_)
);

NAND2_X2 _259_ (
  .A1(_123_),
  .A2(_102_),
  .ZN(_022_)
);

NAND2_X1 _260_ (
  .A1(_021_),
  .A2(_022_),
  .ZN(_023_)
);

NAND2_X1 _261_ (
  .A1(_023_),
  .A2(_117_),
  .ZN(_024_)
);

NAND2_X1 _262_ (
  .A1(_136_),
  .A2(_107_),
  .ZN(_025_)
);

NAND3_X1 _263_ (
  .A1(_024_),
  .A2(_025_),
  .A3(_113_),
  .ZN(_026_)
);

INV_X1 _264_ (
  .A(_009_),
  .ZN(_027_)
);

NAND2_X1 _265_ (
  .A1(_027_),
  .A2(_117_),
  .ZN(_028_)
);

NOR2_X1 _266_ (
  .A1(_119_),
  .A2(_109_),
  .ZN(_029_)
);

NAND2_X1 _267_ (
  .A1(_028_),
  .A2(_029_),
  .ZN(_030_)
);

NAND3_X1 _268_ (
  .A1(_026_),
  .A2(_132_),
  .A3(_030_),
  .ZN(_031_)
);

NAND2_X1 _269_ (
  .A1(_020_),
  .A2(_031_),
  .ZN(_032_)
);

NAND2_X1 _270_ (
  .A1(_144_),
  .A2(\coef[24] ),
  .ZN(_033_)
);

NAND2_X2 _271_ (
  .A1(_032_),
  .A2(_033_),
  .ZN(_002_)
);

NAND3_X2 _272_ (
  .A1(_021_),
  .A2(_022_),
  .A3(_107_),
  .ZN(_034_)
);

NAND2_X1 _273_ (
  .A1(_099_),
  .A2(_101_),
  .ZN(_035_)
);

NAND2_X1 _274_ (
  .A1(_102_),
  .A2(_171_),
  .ZN(_036_)
);

NAND3_X1 _275_ (
  .A1(_035_),
  .A2(_117_),
  .A3(_036_),
  .ZN(_037_)
);

NAND3_X1 _276_ (
  .A1(_034_),
  .A2(_037_),
  .A3(_018_),
  .ZN(_038_)
);

NAND3_X1 _277_ (
  .A1(_152_),
  .A2(_126_),
  .A3(_113_),
  .ZN(_039_)
);

NAND3_X1 _278_ (
  .A1(_038_),
  .A2(_039_),
  .A3(_132_),
  .ZN(_040_)
);

NAND3_X1 _279_ (
  .A1(_118_),
  .A2(_147_),
  .A3(_018_),
  .ZN(_041_)
);

NAND2_X1 _280_ (
  .A1(_099_),
  .A2(_175_),
  .ZN(_042_)
);

NAND2_X1 _281_ (
  .A1(_133_),
  .A2(_102_),
  .ZN(_043_)
);

NAND3_X1 _282_ (
  .A1(_042_),
  .A2(_043_),
  .A3(_107_),
  .ZN(_044_)
);

NAND3_X2 _283_ (
  .A1(_014_),
  .A2(_117_),
  .A3(_015_),
  .ZN(_045_)
);

NAND3_X1 _284_ (
  .A1(_044_),
  .A2(_045_),
  .A3(_109_),
  .ZN(_046_)
);

NAND3_X1 _285_ (
  .A1(_041_),
  .A2(_046_),
  .A3(_097_),
  .ZN(_047_)
);

NAND2_X1 _286_ (
  .A1(_040_),
  .A2(_047_),
  .ZN(_048_)
);

NAND2_X1 _287_ (
  .A1(_048_),
  .A2(_142_),
  .ZN(_049_)
);

NAND2_X1 _288_ (
  .A1(_144_),
  .A2(\coef[10] ),
  .ZN(_050_)
);

NAND2_X1 _289_ (
  .A1(_049_),
  .A2(_050_),
  .ZN(_003_)
);

NAND3_X2 _290_ (
  .A1(_114_),
  .A2(_116_),
  .A3(_107_),
  .ZN(_051_)
);

OAI21_X1 _291_ (
  .A(_051_),
  .B1(_107_),
  .B2(_136_),
  .ZN(_052_)
);

NAND2_X1 _292_ (
  .A1(_052_),
  .A2(_113_),
  .ZN(_053_)
);

NAND2_X1 _293_ (
  .A1(_018_),
  .A2(_165_),
  .ZN(_054_)
);

NAND3_X1 _294_ (
  .A1(_053_),
  .A2(_132_),
  .A3(_054_),
  .ZN(_055_)
);

NAND2_X1 _295_ (
  .A1(_124_),
  .A2(_125_),
  .ZN(_056_)
);

NAND2_X1 _296_ (
  .A1(_056_),
  .A2(_117_),
  .ZN(_057_)
);

NAND3_X1 _297_ (
  .A1(_108_),
  .A2(_057_),
  .A3(_018_),
  .ZN(_058_)
);

OAI21_X1 _298_ (
  .A(_097_),
  .B1(_018_),
  .B2(_165_),
  .ZN(_059_)
);

INV_X1 _299_ (
  .A(_059_),
  .ZN(_060_)
);

AOI21_X1 _300_ (
  .A(_144_),
  .B1(_058_),
  .B2(_060_),
  .ZN(_061_)
);

NAND2_X1 _301_ (
  .A1(_055_),
  .A2(_061_),
  .ZN(_062_)
);

NAND2_X1 _302_ (
  .A1(_144_),
  .A2(\coef[26] ),
  .ZN(_063_)
);

NAND2_X1 _303_ (
  .A1(_062_),
  .A2(_063_),
  .ZN(_004_)
);

NOR2_X1 _304_ (
  .A1(_142_),
  .A2(\coef[13] ),
  .ZN(_064_)
);

NAND3_X1 _305_ (
  .A1(_010_),
  .A2(_018_),
  .A3(_045_),
  .ZN(_065_)
);

NAND3_X1 _306_ (
  .A1(_035_),
  .A2(_107_),
  .A3(_036_),
  .ZN(_066_)
);

NAND2_X1 _307_ (
  .A1(_105_),
  .A2(x[1]),
  .ZN(_067_)
);

NAND2_X1 _308_ (
  .A1(_067_),
  .A2(_109_),
  .ZN(_068_)
);

INV_X1 _309_ (
  .A(_068_),
  .ZN(_069_)
);

AOI21_X1 _310_ (
  .A(_132_),
  .B1(_066_),
  .B2(_069_),
  .ZN(_070_)
);

AOI21_X1 _311_ (
  .A(_144_),
  .B1(_065_),
  .B2(_070_),
  .ZN(_071_)
);

NAND3_X1 _312_ (
  .A1(_028_),
  .A2(_113_),
  .A3(_034_),
  .ZN(_072_)
);

NAND3_X1 _313_ (
  .A1(_042_),
  .A2(_043_),
  .A3(_117_),
  .ZN(_073_)
);

NAND2_X1 _314_ (
  .A1(_107_),
  .A2(_166_),
  .ZN(_074_)
);

NAND3_X1 _315_ (
  .A1(_073_),
  .A2(_018_),
  .A3(_074_),
  .ZN(_075_)
);

NAND3_X1 _316_ (
  .A1(_072_),
  .A2(_075_),
  .A3(_132_),
  .ZN(_076_)
);

AOI21_X1 _317_ (
  .A(_064_),
  .B1(_071_),
  .B2(_076_),
  .ZN(_005_)
);

INV_X1 _318_ (
  .A(_067_),
  .ZN(_077_)
);

OAI21_X1 _319_ (
  .A(_113_),
  .B1(_077_),
  .B2(_138_),
  .ZN(_078_)
);

NAND3_X1 _320_ (
  .A1(_030_),
  .A2(_132_),
  .A3(_078_),
  .ZN(_079_)
);

NAND2_X1 _321_ (
  .A1(_165_),
  .A2(_117_),
  .ZN(_080_)
);

NAND2_X1 _322_ (
  .A1(_107_),
  .A2(x[1]),
  .ZN(_081_)
);

NAND3_X1 _323_ (
  .A1(_080_),
  .A2(_081_),
  .A3(_018_),
  .ZN(_082_)
);

NAND2_X1 _324_ (
  .A1(_013_),
  .A2(_082_),
  .ZN(_083_)
);

NAND3_X1 _325_ (
  .A1(_079_),
  .A2(_083_),
  .A3(_142_),
  .ZN(_084_)
);

NAND2_X1 _326_ (
  .A1(_144_),
  .A2(\coef[28] ),
  .ZN(_085_)
);

NAND2_X1 _327_ (
  .A1(_084_),
  .A2(_085_),
  .ZN(_006_)
);

NAND2_X1 _328_ (
  .A1(_144_),
  .A2(\coef[29] ),
  .ZN(_086_)
);

NAND3_X1 _329_ (
  .A1(_057_),
  .A2(_113_),
  .A3(_081_),
  .ZN(_087_)
);

NAND2_X1 _330_ (
  .A1(_024_),
  .A2(_029_),
  .ZN(_088_)
);

NAND3_X1 _331_ (
  .A1(_087_),
  .A2(_132_),
  .A3(_088_),
  .ZN(_089_)
);

NAND2_X1 _332_ (
  .A1(_089_),
  .A2(_142_),
  .ZN(_090_)
);

NAND3_X1 _333_ (
  .A1(_051_),
  .A2(_018_),
  .A3(_067_),
  .ZN(_091_)
);

NAND2_X1 _334_ (
  .A1(_099_),
  .A2(_117_),
  .ZN(_092_)
);

NAND3_X1 _335_ (
  .A1(_016_),
  .A2(_113_),
  .A3(_092_),
  .ZN(_093_)
);

AOI21_X1 _336_ (
  .A(_132_),
  .B1(_091_),
  .B2(_093_),
  .ZN(_094_)
);

OAI21_X2 _337_ (
  .A(_086_),
  .B1(_090_),
  .B2(_094_),
  .ZN(_007_)
);

NAND3_X1 _338_ (
  .A1(_120_),
  .A2(_142_),
  .A3(_128_),
  .ZN(_095_)
);

INV_X1 _339_ (
  .A(\coef[30] ),
  .ZN(_096_)
);

OAI21_X1 _340_ (
  .A(_095_),
  .B1(_142_),
  .B2(_096_),
  .ZN(_008_)
);

HA_X1 _341_ (
  .A(_165_),
  .B(_166_),
  .CO(_167_),
  .S(_168_)
);

HA_X1 _342_ (
  .A(_165_),
  .B(_166_),
  .CO(_169_),
  .S(_170_)
);

HA_X1 _343_ (
  .A(_165_),
  .B(x[1]),
  .CO(_171_),
  .S(_172_)
);

HA_X1 _344_ (
  .A(_165_),
  .B(x[1]),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _345_ (
  .A(x[0]),
  .B(_166_),
  .CO(_175_),
  .S(_176_)
);

HA_X1 _346_ (
  .A(x[0]),
  .B(_166_),
  .CO(_177_),
  .S(_178_)
);

HA_X1 _347_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_179_),
  .S(_180_)
);

HA_X1 _348_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_181_),
  .S(_182_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_164_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_163_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_162_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_161_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_160_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_159_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_158_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_157_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_156_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$29130e85acc43116076719ea36da8d59b7490cc4\dctu

module \$paramod$4895890460618319d2e2de05b5a45e21ba9e3f8b\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _186_ (
  .A(x[1]),
  .ZN(_169_)
);

INV_X1 _187_ (
  .A(x[0]),
  .ZN(_168_)
);

BUF_X4 _188_ (
  .A(x[2]),
  .Z(_099_)
);

INV_X4 _189_ (
  .A(_099_),
  .ZN(_100_)
);

BUF_X16 _190_ (
  .A(_100_),
  .Z(_101_)
);

NAND2_X2 _191_ (
  .A1(_101_),
  .A2(_170_),
  .ZN(_102_)
);

INV_X1 _192_ (
  .A(_184_),
  .ZN(_103_)
);

BUF_X8 _193_ (
  .A(_099_),
  .Z(_104_)
);

NAND2_X1 _194_ (
  .A1(_103_),
  .A2(_104_),
  .ZN(_105_)
);

BUF_X8 _195_ (
  .A(y[0]),
  .Z(_106_)
);

BUF_X8 _196_ (
  .A(_106_),
  .Z(_107_)
);

NAND3_X1 _197_ (
  .A1(_102_),
  .A2(_105_),
  .A3(_107_),
  .ZN(_108_)
);

NAND2_X4 _198_ (
  .A1(_101_),
  .A2(_178_),
  .ZN(_109_)
);

INV_X1 _199_ (
  .A(_176_),
  .ZN(_110_)
);

NAND2_X2 _200_ (
  .A1(_110_),
  .A2(_104_),
  .ZN(_111_)
);

INV_X8 _201_ (
  .A(_106_),
  .ZN(_112_)
);

BUF_X8 _202_ (
  .A(_112_),
  .Z(_113_)
);

NAND3_X2 _203_ (
  .A1(_109_),
  .A2(_111_),
  .A3(_113_),
  .ZN(_114_)
);

BUF_X2 _204_ (
  .A(y[1]),
  .Z(_115_)
);

INV_X1 _205_ (
  .A(_115_),
  .ZN(_116_)
);

NAND3_X1 _206_ (
  .A1(_108_),
  .A2(_114_),
  .A3(_116_),
  .ZN(_117_)
);

NAND2_X1 _207_ (
  .A1(_100_),
  .A2(_182_),
  .ZN(_118_)
);

INV_X1 _208_ (
  .A(_172_),
  .ZN(_119_)
);

NAND2_X1 _209_ (
  .A1(_119_),
  .A2(_099_),
  .ZN(_120_)
);

NAND3_X1 _210_ (
  .A1(_118_),
  .A2(_120_),
  .A3(_106_),
  .ZN(_121_)
);

NAND2_X4 _211_ (
  .A1(_101_),
  .A2(_174_),
  .ZN(_122_)
);

INV_X1 _212_ (
  .A(_180_),
  .ZN(_123_)
);

NAND2_X1 _213_ (
  .A1(_123_),
  .A2(_099_),
  .ZN(_124_)
);

NAND3_X2 _214_ (
  .A1(_122_),
  .A2(_124_),
  .A3(_112_),
  .ZN(_125_)
);

BUF_X2 _215_ (
  .A(_115_),
  .Z(_126_)
);

NAND3_X1 _216_ (
  .A1(_121_),
  .A2(_125_),
  .A3(_126_),
  .ZN(_127_)
);

BUF_X2 _217_ (
  .A(y[2]),
  .Z(_128_)
);

INV_X1 _218_ (
  .A(_128_),
  .ZN(_129_)
);

NAND3_X1 _219_ (
  .A1(_117_),
  .A2(_127_),
  .A3(_129_),
  .ZN(_130_)
);

NAND2_X4 _220_ (
  .A1(_101_),
  .A2(_110_),
  .ZN(_131_)
);

NAND2_X4 _221_ (
  .A1(_104_),
  .A2(_178_),
  .ZN(_132_)
);

NAND3_X4 _222_ (
  .A1(_131_),
  .A2(_106_),
  .A3(_132_),
  .ZN(_133_)
);

NAND2_X4 _223_ (
  .A1(_101_),
  .A2(_103_),
  .ZN(_134_)
);

NAND2_X2 _224_ (
  .A1(_104_),
  .A2(_170_),
  .ZN(_135_)
);

NAND3_X2 _225_ (
  .A1(_134_),
  .A2(_113_),
  .A3(_135_),
  .ZN(_136_)
);

NAND3_X1 _226_ (
  .A1(_133_),
  .A2(_136_),
  .A3(_116_),
  .ZN(_137_)
);

NAND2_X4 _227_ (
  .A1(_101_),
  .A2(_123_),
  .ZN(_138_)
);

NAND2_X2 _228_ (
  .A1(_104_),
  .A2(_174_),
  .ZN(_139_)
);

NAND3_X2 _229_ (
  .A1(_138_),
  .A2(_106_),
  .A3(_139_),
  .ZN(_140_)
);

NAND2_X2 _230_ (
  .A1(_101_),
  .A2(_119_),
  .ZN(_141_)
);

NAND2_X1 _231_ (
  .A1(_104_),
  .A2(_182_),
  .ZN(_142_)
);

NAND3_X1 _232_ (
  .A1(_141_),
  .A2(_113_),
  .A3(_142_),
  .ZN(_143_)
);

NAND3_X1 _233_ (
  .A1(_140_),
  .A2(_143_),
  .A3(_115_),
  .ZN(_144_)
);

NAND3_X1 _234_ (
  .A1(_137_),
  .A2(_144_),
  .A3(_128_),
  .ZN(_145_)
);

NAND2_X1 _235_ (
  .A1(_130_),
  .A2(_145_),
  .ZN(_146_)
);

BUF_X2 _236_ (
  .A(ena),
  .Z(_147_)
);

NAND2_X1 _237_ (
  .A1(_146_),
  .A2(_147_),
  .ZN(_148_)
);

INV_X1 _238_ (
  .A(ena),
  .ZN(_149_)
);

NAND2_X1 _239_ (
  .A1(_149_),
  .A2(\coef[10] ),
  .ZN(_150_)
);

NAND2_X1 _240_ (
  .A1(_148_),
  .A2(_150_),
  .ZN(_000_)
);

NAND2_X1 _241_ (
  .A1(_141_),
  .A2(_142_),
  .ZN(_151_)
);

NAND2_X1 _242_ (
  .A1(_151_),
  .A2(_107_),
  .ZN(_152_)
);

INV_X1 _243_ (
  .A(_171_),
  .ZN(_153_)
);

NAND2_X4 _244_ (
  .A1(_101_),
  .A2(_153_),
  .ZN(_154_)
);

NAND2_X1 _245_ (
  .A1(_099_),
  .A2(_171_),
  .ZN(_155_)
);

NAND2_X4 _246_ (
  .A1(_154_),
  .A2(_155_),
  .ZN(_156_)
);

NAND2_X4 _247_ (
  .A1(_156_),
  .A2(_113_),
  .ZN(_157_)
);

BUF_X4 _248_ (
  .A(_116_),
  .Z(_158_)
);

NAND3_X1 _249_ (
  .A1(_152_),
  .A2(_157_),
  .A3(_158_),
  .ZN(_009_)
);

NAND2_X2 _250_ (
  .A1(_107_),
  .A2(x[1]),
  .ZN(_010_)
);

NAND2_X1 _251_ (
  .A1(_114_),
  .A2(_010_),
  .ZN(_011_)
);

NAND2_X1 _252_ (
  .A1(_011_),
  .A2(_126_),
  .ZN(_012_)
);

NAND3_X1 _253_ (
  .A1(_009_),
  .A2(_012_),
  .A3(_129_),
  .ZN(_013_)
);

NAND2_X1 _254_ (
  .A1(_102_),
  .A2(_105_),
  .ZN(_014_)
);

NAND2_X1 _255_ (
  .A1(_014_),
  .A2(_113_),
  .ZN(_015_)
);

NAND3_X2 _256_ (
  .A1(_154_),
  .A2(_107_),
  .A3(_155_),
  .ZN(_016_)
);

NAND3_X1 _257_ (
  .A1(_015_),
  .A2(_016_),
  .A3(_126_),
  .ZN(_017_)
);

NAND2_X2 _258_ (
  .A1(_113_),
  .A2(_169_),
  .ZN(_018_)
);

NAND2_X1 _259_ (
  .A1(_140_),
  .A2(_018_),
  .ZN(_019_)
);

NAND2_X1 _260_ (
  .A1(_019_),
  .A2(_158_),
  .ZN(_020_)
);

NAND3_X1 _261_ (
  .A1(_017_),
  .A2(_020_),
  .A3(_128_),
  .ZN(_021_)
);

NAND3_X1 _262_ (
  .A1(_013_),
  .A2(_021_),
  .A3(_147_),
  .ZN(_022_)
);

NAND2_X1 _263_ (
  .A1(_149_),
  .A2(\coef[13] ),
  .ZN(_023_)
);

NAND2_X1 _264_ (
  .A1(_022_),
  .A2(_023_),
  .ZN(_001_)
);

INV_X1 _265_ (
  .A(_133_),
  .ZN(_024_)
);

NOR2_X2 _266_ (
  .A1(_106_),
  .A2(x[0]),
  .ZN(_025_)
);

OAI21_X1 _267_ (
  .A(_158_),
  .B1(_024_),
  .B2(_025_),
  .ZN(_026_)
);

NAND2_X1 _268_ (
  .A1(_118_),
  .A2(_120_),
  .ZN(_027_)
);

NAND2_X1 _269_ (
  .A1(_027_),
  .A2(_113_),
  .ZN(_028_)
);

OAI21_X2 _270_ (
  .A(_115_),
  .B1(_112_),
  .B2(_104_),
  .ZN(_029_)
);

INV_X1 _271_ (
  .A(_029_),
  .ZN(_030_)
);

AOI21_X1 _272_ (
  .A(_128_),
  .B1(_028_),
  .B2(_030_),
  .ZN(_031_)
);

AOI21_X2 _273_ (
  .A(_149_),
  .B1(_026_),
  .B2(_031_),
  .ZN(_032_)
);

NAND2_X2 _274_ (
  .A1(_106_),
  .A2(x[0]),
  .ZN(_033_)
);

NAND2_X1 _275_ (
  .A1(_125_),
  .A2(_033_),
  .ZN(_034_)
);

NAND2_X1 _276_ (
  .A1(_034_),
  .A2(_126_),
  .ZN(_035_)
);

NAND2_X4 _277_ (
  .A1(_134_),
  .A2(_135_),
  .ZN(_036_)
);

NAND2_X2 _278_ (
  .A1(_036_),
  .A2(_107_),
  .ZN(_037_)
);

NOR2_X4 _279_ (
  .A1(_101_),
  .A2(_106_),
  .ZN(_038_)
);

INV_X2 _280_ (
  .A(_038_),
  .ZN(_039_)
);

NAND3_X1 _281_ (
  .A1(_037_),
  .A2(_158_),
  .A3(_039_),
  .ZN(_040_)
);

NAND3_X1 _282_ (
  .A1(_035_),
  .A2(_040_),
  .A3(_128_),
  .ZN(_041_)
);

NAND2_X2 _283_ (
  .A1(_032_),
  .A2(_041_),
  .ZN(_042_)
);

NAND2_X1 _284_ (
  .A1(_149_),
  .A2(\coef[21] ),
  .ZN(_043_)
);

NAND2_X2 _285_ (
  .A1(_042_),
  .A2(_043_),
  .ZN(_002_)
);

NAND2_X1 _286_ (
  .A1(_039_),
  .A2(_116_),
  .ZN(_044_)
);

OAI21_X1 _287_ (
  .A(_044_),
  .B1(_158_),
  .B2(_025_),
  .ZN(_045_)
);

NAND3_X1 _288_ (
  .A1(_045_),
  .A2(_128_),
  .A3(_121_),
  .ZN(_046_)
);

INV_X1 _289_ (
  .A(_033_),
  .ZN(_047_)
);

OAI21_X1 _290_ (
  .A(_029_),
  .B1(_126_),
  .B2(_047_),
  .ZN(_048_)
);

NAND3_X1 _291_ (
  .A1(_048_),
  .A2(_129_),
  .A3(_136_),
  .ZN(_049_)
);

NAND3_X1 _292_ (
  .A1(_046_),
  .A2(_049_),
  .A3(_147_),
  .ZN(_050_)
);

INV_X1 _293_ (
  .A(\coef[23] ),
  .ZN(_051_)
);

OAI21_X1 _294_ (
  .A(_050_),
  .B1(_147_),
  .B2(_051_),
  .ZN(_003_)
);

NAND2_X2 _295_ (
  .A1(_138_),
  .A2(_139_),
  .ZN(_052_)
);

NAND2_X2 _296_ (
  .A1(_052_),
  .A2(_113_),
  .ZN(_053_)
);

NAND2_X1 _297_ (
  .A1(_027_),
  .A2(_107_),
  .ZN(_054_)
);

NAND3_X1 _298_ (
  .A1(_053_),
  .A2(_054_),
  .A3(_158_),
  .ZN(_055_)
);

NAND2_X1 _299_ (
  .A1(_033_),
  .A2(_115_),
  .ZN(_056_)
);

INV_X1 _300_ (
  .A(_056_),
  .ZN(_057_)
);

AOI21_X2 _301_ (
  .A(_129_),
  .B1(_057_),
  .B2(_018_),
  .ZN(_058_)
);

NAND2_X1 _302_ (
  .A1(_055_),
  .A2(_058_),
  .ZN(_059_)
);

NAND2_X2 _303_ (
  .A1(_109_),
  .A2(_111_),
  .ZN(_060_)
);

NAND2_X2 _304_ (
  .A1(_060_),
  .A2(_107_),
  .ZN(_061_)
);

NAND2_X2 _305_ (
  .A1(_036_),
  .A2(_113_),
  .ZN(_062_)
);

NAND3_X1 _306_ (
  .A1(_061_),
  .A2(_062_),
  .A3(_126_),
  .ZN(_063_)
);

NOR2_X2 _307_ (
  .A1(_025_),
  .A2(_115_),
  .ZN(_064_)
);

AOI21_X2 _308_ (
  .A(_128_),
  .B1(_064_),
  .B2(_010_),
  .ZN(_065_)
);

NAND2_X1 _309_ (
  .A1(_063_),
  .A2(_065_),
  .ZN(_066_)
);

NAND3_X1 _310_ (
  .A1(_059_),
  .A2(_066_),
  .A3(_147_),
  .ZN(_067_)
);

INV_X1 _311_ (
  .A(\coef[24] ),
  .ZN(_068_)
);

OAI21_X1 _312_ (
  .A(_067_),
  .B1(_147_),
  .B2(_068_),
  .ZN(_004_)
);

NAND2_X4 _313_ (
  .A1(_131_),
  .A2(_132_),
  .ZN(_069_)
);

NAND2_X4 _314_ (
  .A1(_069_),
  .A2(_113_),
  .ZN(_070_)
);

NAND3_X2 _315_ (
  .A1(_037_),
  .A2(_070_),
  .A3(_126_),
  .ZN(_071_)
);

AOI21_X1 _316_ (
  .A(_128_),
  .B1(_158_),
  .B2(_104_),
  .ZN(_072_)
);

AOI21_X2 _317_ (
  .A(_149_),
  .B1(_071_),
  .B2(_072_),
  .ZN(_073_)
);

NAND2_X2 _318_ (
  .A1(_122_),
  .A2(_124_),
  .ZN(_074_)
);

NAND2_X2 _319_ (
  .A1(_074_),
  .A2(_107_),
  .ZN(_075_)
);

NAND3_X1 _320_ (
  .A1(_028_),
  .A2(_075_),
  .A3(_158_),
  .ZN(_076_)
);

NAND2_X1 _321_ (
  .A1(_101_),
  .A2(_126_),
  .ZN(_077_)
);

NAND3_X1 _322_ (
  .A1(_076_),
  .A2(_128_),
  .A3(_077_),
  .ZN(_078_)
);

NAND2_X1 _323_ (
  .A1(_073_),
  .A2(_078_),
  .ZN(_079_)
);

NAND2_X1 _324_ (
  .A1(_149_),
  .A2(\coef[26] ),
  .ZN(_080_)
);

NAND2_X1 _325_ (
  .A1(_079_),
  .A2(_080_),
  .ZN(_005_)
);

INV_X1 _326_ (
  .A(_016_),
  .ZN(_081_)
);

OAI21_X1 _327_ (
  .A(_126_),
  .B1(_104_),
  .B2(_107_),
  .ZN(_082_)
);

OAI21_X1 _328_ (
  .A(_065_),
  .B1(_081_),
  .B2(_082_),
  .ZN(_083_)
);

NAND2_X1 _329_ (
  .A1(_104_),
  .A2(_107_),
  .ZN(_084_)
);

NAND3_X1 _330_ (
  .A1(_157_),
  .A2(_158_),
  .A3(_084_),
  .ZN(_085_)
);

NAND2_X1 _331_ (
  .A1(_085_),
  .A2(_058_),
  .ZN(_086_)
);

NAND3_X1 _332_ (
  .A1(_083_),
  .A2(_147_),
  .A3(_086_),
  .ZN(_087_)
);

INV_X1 _333_ (
  .A(\coef[28] ),
  .ZN(_088_)
);

OAI21_X1 _334_ (
  .A(_087_),
  .B1(_147_),
  .B2(_088_),
  .ZN(_006_)
);

AOI21_X1 _335_ (
  .A(_128_),
  .B1(_061_),
  .B2(_064_),
  .ZN(_089_)
);

NAND3_X1 _336_ (
  .A1(_157_),
  .A2(_075_),
  .A3(_126_),
  .ZN(_090_)
);

NAND2_X1 _337_ (
  .A1(_089_),
  .A2(_090_),
  .ZN(_091_)
);

AOI21_X1 _338_ (
  .A(_129_),
  .B1(_053_),
  .B2(_057_),
  .ZN(_092_)
);

NAND3_X1 _339_ (
  .A1(_070_),
  .A2(_016_),
  .A3(_158_),
  .ZN(_093_)
);

NAND2_X1 _340_ (
  .A1(_092_),
  .A2(_093_),
  .ZN(_094_)
);

NAND3_X1 _341_ (
  .A1(_091_),
  .A2(_094_),
  .A3(_147_),
  .ZN(_095_)
);

NAND2_X1 _342_ (
  .A1(_149_),
  .A2(\coef[29] ),
  .ZN(_096_)
);

NAND2_X1 _343_ (
  .A1(_095_),
  .A2(_096_),
  .ZN(_007_)
);

NAND2_X1 _344_ (
  .A1(_149_),
  .A2(\coef[30] ),
  .ZN(_097_)
);

NAND2_X1 _345_ (
  .A1(_033_),
  .A2(_147_),
  .ZN(_098_)
);

OAI21_X1 _346_ (
  .A(_097_),
  .B1(_098_),
  .B2(_025_),
  .ZN(_008_)
);

HA_X1 _347_ (
  .A(_168_),
  .B(_169_),
  .CO(_170_),
  .S(_171_)
);

HA_X1 _348_ (
  .A(_168_),
  .B(_169_),
  .CO(_172_),
  .S(_173_)
);

HA_X1 _349_ (
  .A(_168_),
  .B(x[1]),
  .CO(_174_),
  .S(_175_)
);

HA_X1 _350_ (
  .A(_168_),
  .B(x[1]),
  .CO(_176_),
  .S(_177_)
);

HA_X1 _351_ (
  .A(x[0]),
  .B(_169_),
  .CO(_178_),
  .S(_179_)
);

HA_X1 _352_ (
  .A(x[0]),
  .B(_169_),
  .CO(_180_),
  .S(_181_)
);

HA_X1 _353_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_182_),
  .S(_183_)
);

HA_X1 _354_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_184_),
  .S(_185_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_165_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_164_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_163_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_167_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_162_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_166_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_161_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_160_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_159_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$4895890460618319d2e2de05b5a45e21ba9e3f8b\dctu

module \$paramod$4dc5718e86f31fe555f7d39cf5ab7078c09f577a\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _189_ (
  .A(x[1]),
  .ZN(_172_)
);

INV_X1 _190_ (
  .A(x[0]),
  .ZN(_171_)
);

BUF_X1 _191_ (
  .A(ena),
  .Z(_103_)
);

NOR2_X1 _192_ (
  .A1(\coef[21] ),
  .A2(_103_),
  .ZN(_104_)
);

BUF_X4 _193_ (
  .A(y[1]),
  .Z(_105_)
);

INV_X4 _194_ (
  .A(_105_),
  .ZN(_106_)
);

BUF_X2 _195_ (
  .A(y[2]),
  .Z(_107_)
);

NOR2_X4 _196_ (
  .A1(_106_),
  .A2(_107_),
  .ZN(_108_)
);

INV_X1 _197_ (
  .A(_108_),
  .ZN(_109_)
);

INV_X2 _198_ (
  .A(x[2]),
  .ZN(_110_)
);

INV_X1 _199_ (
  .A(_175_),
  .ZN(_111_)
);

NAND2_X1 _200_ (
  .A1(_110_),
  .A2(_111_),
  .ZN(_112_)
);

BUF_X4 _201_ (
  .A(x[2]),
  .Z(_113_)
);

NAND2_X4 _202_ (
  .A1(_113_),
  .A2(_185_),
  .ZN(_114_)
);

NAND2_X4 _203_ (
  .A1(_112_),
  .A2(_114_),
  .ZN(_115_)
);

BUF_X4 _204_ (
  .A(y[0]),
  .Z(_116_)
);

INV_X4 _205_ (
  .A(_116_),
  .ZN(_117_)
);

BUF_X8 _206_ (
  .A(_117_),
  .Z(_118_)
);

AOI21_X4 _207_ (
  .A(_109_),
  .B1(_115_),
  .B2(_118_),
  .ZN(_119_)
);

INV_X1 _208_ (
  .A(_179_),
  .ZN(_120_)
);

NAND2_X1 _209_ (
  .A1(_110_),
  .A2(_120_),
  .ZN(_121_)
);

NAND2_X1 _210_ (
  .A1(_113_),
  .A2(_181_),
  .ZN(_122_)
);

NAND2_X1 _211_ (
  .A1(_121_),
  .A2(_122_),
  .ZN(_123_)
);

BUF_X4 _212_ (
  .A(_116_),
  .Z(_124_)
);

NAND2_X1 _213_ (
  .A1(_123_),
  .A2(_124_),
  .ZN(_125_)
);

NAND2_X1 _214_ (
  .A1(_119_),
  .A2(_125_),
  .ZN(_126_)
);

INV_X1 _215_ (
  .A(_173_),
  .ZN(_127_)
);

NAND2_X1 _216_ (
  .A1(_110_),
  .A2(_127_),
  .ZN(_128_)
);

NAND2_X4 _217_ (
  .A1(_113_),
  .A2(_187_),
  .ZN(_129_)
);

NAND3_X2 _218_ (
  .A1(_128_),
  .A2(_118_),
  .A3(_129_),
  .ZN(_130_)
);

INV_X1 _219_ (
  .A(_177_),
  .ZN(_131_)
);

NAND2_X1 _220_ (
  .A1(_110_),
  .A2(_131_),
  .ZN(_132_)
);

NAND2_X1 _221_ (
  .A1(_113_),
  .A2(_183_),
  .ZN(_133_)
);

NAND3_X1 _222_ (
  .A1(_132_),
  .A2(_124_),
  .A3(_133_),
  .ZN(_134_)
);

NAND2_X1 _223_ (
  .A1(_105_),
  .A2(_107_),
  .ZN(_135_)
);

INV_X1 _224_ (
  .A(_135_),
  .ZN(_136_)
);

NAND3_X1 _225_ (
  .A1(_130_),
  .A2(_134_),
  .A3(_136_),
  .ZN(_137_)
);

NAND2_X1 _226_ (
  .A1(_126_),
  .A2(_137_),
  .ZN(_138_)
);

NAND2_X2 _227_ (
  .A1(_106_),
  .A2(_107_),
  .ZN(_139_)
);

INV_X1 _228_ (
  .A(_115_),
  .ZN(_140_)
);

NAND2_X1 _229_ (
  .A1(_140_),
  .A2(_124_),
  .ZN(_141_)
);

NAND3_X1 _230_ (
  .A1(_121_),
  .A2(_118_),
  .A3(_122_),
  .ZN(_142_)
);

AOI21_X1 _231_ (
  .A(_139_),
  .B1(_141_),
  .B2(_142_),
  .ZN(_143_)
);

NOR2_X2 _232_ (
  .A1(_138_),
  .A2(_143_),
  .ZN(_144_)
);

INV_X1 _233_ (
  .A(_103_),
  .ZN(_145_)
);

NAND2_X1 _234_ (
  .A1(_128_),
  .A2(_129_),
  .ZN(_146_)
);

NAND2_X1 _235_ (
  .A1(_146_),
  .A2(_116_),
  .ZN(_147_)
);

NAND2_X2 _236_ (
  .A1(_132_),
  .A2(_133_),
  .ZN(_148_)
);

INV_X1 _237_ (
  .A(_148_),
  .ZN(_149_)
);

OAI21_X1 _238_ (
  .A(_147_),
  .B1(_149_),
  .B2(_124_),
  .ZN(_150_)
);

NOR2_X1 _239_ (
  .A1(_105_),
  .A2(_107_),
  .ZN(_151_)
);

AOI21_X1 _240_ (
  .A(_145_),
  .B1(_150_),
  .B2(_151_),
  .ZN(_152_)
);

AOI21_X2 _241_ (
  .A(_104_),
  .B1(_144_),
  .B2(_152_),
  .ZN(_000_)
);

NAND2_X1 _242_ (
  .A1(_110_),
  .A2(_181_),
  .ZN(_153_)
);

NAND2_X1 _243_ (
  .A1(_120_),
  .A2(_113_),
  .ZN(_154_)
);

NAND3_X1 _244_ (
  .A1(_153_),
  .A2(_154_),
  .A3(_118_),
  .ZN(_155_)
);

INV_X1 _245_ (
  .A(_183_),
  .ZN(_156_)
);

NAND2_X1 _246_ (
  .A1(_110_),
  .A2(_156_),
  .ZN(_157_)
);

NAND2_X1 _247_ (
  .A1(_113_),
  .A2(_177_),
  .ZN(_158_)
);

NAND3_X1 _248_ (
  .A1(_157_),
  .A2(_116_),
  .A3(_158_),
  .ZN(_159_)
);

NAND3_X1 _249_ (
  .A1(_155_),
  .A2(_159_),
  .A3(_107_),
  .ZN(_160_)
);

NAND3_X1 _250_ (
  .A1(_153_),
  .A2(_154_),
  .A3(_116_),
  .ZN(_010_)
);

NAND3_X1 _251_ (
  .A1(_157_),
  .A2(_118_),
  .A3(_158_),
  .ZN(_011_)
);

INV_X1 _252_ (
  .A(_107_),
  .ZN(_012_)
);

NAND3_X1 _253_ (
  .A1(_010_),
  .A2(_011_),
  .A3(_012_),
  .ZN(_013_)
);

BUF_X1 _254_ (
  .A(_103_),
  .Z(_014_)
);

NAND3_X1 _255_ (
  .A1(_160_),
  .A2(_013_),
  .A3(_014_),
  .ZN(_015_)
);

INV_X1 _256_ (
  .A(\coef[22] ),
  .ZN(_016_)
);

OAI21_X1 _257_ (
  .A(_015_),
  .B1(_014_),
  .B2(_016_),
  .ZN(_001_)
);

NOR2_X1 _258_ (
  .A1(_014_),
  .A2(\coef[23] ),
  .ZN(_017_)
);

NAND2_X1 _259_ (
  .A1(_113_),
  .A2(_116_),
  .ZN(_018_)
);

NAND2_X1 _260_ (
  .A1(_018_),
  .A2(_105_),
  .ZN(_019_)
);

INV_X1 _261_ (
  .A(_019_),
  .ZN(_020_)
);

OAI21_X1 _262_ (
  .A(_020_),
  .B1(_148_),
  .B2(_124_),
  .ZN(_021_)
);

NOR2_X1 _263_ (
  .A1(_113_),
  .A2(_116_),
  .ZN(_022_)
);

NOR2_X1 _264_ (
  .A1(_022_),
  .A2(_105_),
  .ZN(_023_)
);

NAND2_X1 _265_ (
  .A1(_125_),
  .A2(_023_),
  .ZN(_024_)
);

NAND2_X1 _266_ (
  .A1(_021_),
  .A2(_024_),
  .ZN(_025_)
);

AOI21_X1 _267_ (
  .A(_145_),
  .B1(_025_),
  .B2(_012_),
  .ZN(_026_)
);

AOI21_X1 _268_ (
  .A(_012_),
  .B1(_142_),
  .B2(_020_),
  .ZN(_027_)
);

OAI21_X1 _269_ (
  .A(_023_),
  .B1(_149_),
  .B2(_118_),
  .ZN(_028_)
);

NAND2_X1 _270_ (
  .A1(_027_),
  .A2(_028_),
  .ZN(_029_)
);

AOI21_X1 _271_ (
  .A(_017_),
  .B1(_026_),
  .B2(_029_),
  .ZN(_002_)
);

INV_X1 _272_ (
  .A(_018_),
  .ZN(_030_)
);

NOR2_X1 _273_ (
  .A1(_030_),
  .A2(_022_),
  .ZN(_031_)
);

XNOR2_X1 _274_ (
  .A(_107_),
  .B(_174_),
  .ZN(_032_)
);

OR2_X1 _275_ (
  .A1(_031_),
  .A2(_032_),
  .ZN(_033_)
);

NAND2_X1 _276_ (
  .A1(_031_),
  .A2(_032_),
  .ZN(_034_)
);

NAND3_X1 _277_ (
  .A1(_033_),
  .A2(_034_),
  .A3(_014_),
  .ZN(_035_)
);

INV_X1 _278_ (
  .A(\coef[24] ),
  .ZN(_036_)
);

OAI21_X1 _279_ (
  .A(_035_),
  .B1(_014_),
  .B2(_036_),
  .ZN(_003_)
);

AOI21_X1 _280_ (
  .A(_139_),
  .B1(x[1]),
  .B2(_118_),
  .ZN(_037_)
);

NAND2_X4 _281_ (
  .A1(_115_),
  .A2(_124_),
  .ZN(_038_)
);

AOI21_X1 _282_ (
  .A(_145_),
  .B1(_037_),
  .B2(_038_),
  .ZN(_039_)
);

INV_X1 _283_ (
  .A(_146_),
  .ZN(_040_)
);

NAND2_X1 _284_ (
  .A1(_040_),
  .A2(_124_),
  .ZN(_041_)
);

NOR2_X1 _285_ (
  .A1(_116_),
  .A2(x[1]),
  .ZN(_042_)
);

INV_X1 _286_ (
  .A(_042_),
  .ZN(_043_)
);

NAND3_X1 _287_ (
  .A1(_041_),
  .A2(_151_),
  .A3(_043_),
  .ZN(_044_)
);

NAND2_X1 _288_ (
  .A1(_039_),
  .A2(_044_),
  .ZN(_045_)
);

NAND2_X1 _289_ (
  .A1(_124_),
  .A2(x[1]),
  .ZN(_046_)
);

NAND2_X1 _290_ (
  .A1(_119_),
  .A2(_046_),
  .ZN(_047_)
);

NAND2_X1 _291_ (
  .A1(_172_),
  .A2(_124_),
  .ZN(_048_)
);

NAND3_X1 _292_ (
  .A1(_130_),
  .A2(_136_),
  .A3(_048_),
  .ZN(_049_)
);

NAND2_X1 _293_ (
  .A1(_047_),
  .A2(_049_),
  .ZN(_050_)
);

NOR2_X1 _294_ (
  .A1(_045_),
  .A2(_050_),
  .ZN(_051_)
);

NOR2_X1 _295_ (
  .A1(_014_),
  .A2(\coef[25] ),
  .ZN(_052_)
);

NOR2_X2 _296_ (
  .A1(_051_),
  .A2(_052_),
  .ZN(_004_)
);

NOR2_X1 _297_ (
  .A1(_014_),
  .A2(\coef[26] ),
  .ZN(_053_)
);

AOI21_X2 _298_ (
  .A(_106_),
  .B1(_171_),
  .B2(_118_),
  .ZN(_054_)
);

NAND2_X1 _299_ (
  .A1(_038_),
  .A2(_054_),
  .ZN(_055_)
);

OAI21_X1 _300_ (
  .A(_106_),
  .B1(_117_),
  .B2(_171_),
  .ZN(_056_)
);

INV_X1 _301_ (
  .A(_056_),
  .ZN(_057_)
);

NAND2_X1 _302_ (
  .A1(_130_),
  .A2(_057_),
  .ZN(_058_)
);

NAND2_X1 _303_ (
  .A1(_055_),
  .A2(_058_),
  .ZN(_059_)
);

AOI21_X1 _304_ (
  .A(_145_),
  .B1(_059_),
  .B2(_012_),
  .ZN(_060_)
);

AOI21_X1 _305_ (
  .A(_012_),
  .B1(_147_),
  .B2(_054_),
  .ZN(_061_)
);

OAI21_X1 _306_ (
  .A(_057_),
  .B1(_124_),
  .B2(_115_),
  .ZN(_062_)
);

NAND2_X1 _307_ (
  .A1(_061_),
  .A2(_062_),
  .ZN(_063_)
);

AOI21_X2 _308_ (
  .A(_053_),
  .B1(_060_),
  .B2(_063_),
  .ZN(_005_)
);

NAND2_X1 _309_ (
  .A1(_110_),
  .A2(_185_),
  .ZN(_064_)
);

NAND2_X1 _310_ (
  .A1(_111_),
  .A2(_113_),
  .ZN(_065_)
);

NAND3_X1 _311_ (
  .A1(_064_),
  .A2(_065_),
  .A3(_116_),
  .ZN(_066_)
);

NAND2_X1 _312_ (
  .A1(_155_),
  .A2(_066_),
  .ZN(_067_)
);

NAND2_X1 _313_ (
  .A1(_067_),
  .A2(_108_),
  .ZN(_068_)
);

NAND3_X1 _314_ (
  .A1(_064_),
  .A2(_065_),
  .A3(_118_),
  .ZN(_069_)
);

NAND2_X1 _315_ (
  .A1(_010_),
  .A2(_069_),
  .ZN(_070_)
);

INV_X1 _316_ (
  .A(_139_),
  .ZN(_071_)
);

NAND2_X1 _317_ (
  .A1(_070_),
  .A2(_071_),
  .ZN(_072_)
);

INV_X1 _318_ (
  .A(_187_),
  .ZN(_073_)
);

NAND2_X1 _319_ (
  .A1(_110_),
  .A2(_073_),
  .ZN(_074_)
);

NAND2_X1 _320_ (
  .A1(_113_),
  .A2(_173_),
  .ZN(_075_)
);

NAND3_X1 _321_ (
  .A1(_074_),
  .A2(_116_),
  .A3(_075_),
  .ZN(_076_)
);

NAND2_X1 _322_ (
  .A1(_011_),
  .A2(_076_),
  .ZN(_077_)
);

NAND2_X1 _323_ (
  .A1(_077_),
  .A2(_136_),
  .ZN(_078_)
);

NAND3_X1 _324_ (
  .A1(_068_),
  .A2(_072_),
  .A3(_078_),
  .ZN(_079_)
);

NAND3_X1 _325_ (
  .A1(_074_),
  .A2(_118_),
  .A3(_075_),
  .ZN(_080_)
);

NAND2_X1 _326_ (
  .A1(_159_),
  .A2(_080_),
  .ZN(_081_)
);

NAND2_X1 _327_ (
  .A1(_081_),
  .A2(_151_),
  .ZN(_082_)
);

NAND2_X1 _328_ (
  .A1(_082_),
  .A2(_103_),
  .ZN(_083_)
);

NOR2_X1 _329_ (
  .A1(_079_),
  .A2(_083_),
  .ZN(_084_)
);

NOR2_X1 _330_ (
  .A1(_014_),
  .A2(\coef[27] ),
  .ZN(_085_)
);

NOR2_X1 _331_ (
  .A1(_084_),
  .A2(_085_),
  .ZN(_006_)
);

NOR2_X1 _332_ (
  .A1(_103_),
  .A2(\coef[28] ),
  .ZN(_086_)
);

NOR2_X2 _333_ (
  .A1(_071_),
  .A2(_108_),
  .ZN(_087_)
);

AOI21_X1 _334_ (
  .A(_145_),
  .B1(_087_),
  .B2(_148_),
  .ZN(_088_)
);

OR2_X1 _335_ (
  .A1(_087_),
  .A2(_123_),
  .ZN(_089_)
);

AOI21_X1 _336_ (
  .A(_086_),
  .B1(_088_),
  .B2(_089_),
  .ZN(_007_)
);

NOR2_X1 _337_ (
  .A1(_042_),
  .A2(_139_),
  .ZN(_090_)
);

AOI21_X1 _338_ (
  .A(_145_),
  .B1(_038_),
  .B2(_090_),
  .ZN(_091_)
);

NAND2_X1 _339_ (
  .A1(_147_),
  .A2(_043_),
  .ZN(_092_)
);

NAND2_X1 _340_ (
  .A1(_092_),
  .A2(_151_),
  .ZN(_093_)
);

NAND2_X1 _341_ (
  .A1(_091_),
  .A2(_093_),
  .ZN(_094_)
);

NAND2_X1 _342_ (
  .A1(_119_),
  .A2(_048_),
  .ZN(_095_)
);

NAND3_X1 _343_ (
  .A1(_130_),
  .A2(_136_),
  .A3(_046_),
  .ZN(_096_)
);

NAND2_X1 _344_ (
  .A1(_095_),
  .A2(_096_),
  .ZN(_097_)
);

NOR2_X1 _345_ (
  .A1(_094_),
  .A2(_097_),
  .ZN(_098_)
);

NOR2_X1 _346_ (
  .A1(_014_),
  .A2(\coef[15] ),
  .ZN(_099_)
);

NOR2_X2 _347_ (
  .A1(_098_),
  .A2(_099_),
  .ZN(_008_)
);

AOI21_X1 _348_ (
  .A(_145_),
  .B1(_087_),
  .B2(_040_),
  .ZN(_100_)
);

OAI21_X1 _349_ (
  .A(_100_),
  .B1(_140_),
  .B2(_087_),
  .ZN(_101_)
);

INV_X1 _350_ (
  .A(\coef[30] ),
  .ZN(_102_)
);

OAI21_X1 _351_ (
  .A(_101_),
  .B1(_014_),
  .B2(_102_),
  .ZN(_009_)
);

HA_X1 _352_ (
  .A(_171_),
  .B(_172_),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _353_ (
  .A(_171_),
  .B(_172_),
  .CO(_175_),
  .S(_176_)
);

HA_X1 _354_ (
  .A(_171_),
  .B(x[1]),
  .CO(_177_),
  .S(_178_)
);

HA_X1 _355_ (
  .A(_171_),
  .B(x[1]),
  .CO(_179_),
  .S(_180_)
);

HA_X1 _356_ (
  .A(x[0]),
  .B(_172_),
  .CO(_181_),
  .S(_182_)
);

HA_X1 _357_ (
  .A(x[0]),
  .B(_172_),
  .CO(_183_),
  .S(_184_)
);

HA_X1 _358_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_185_),
  .S(_186_)
);

HA_X1 _359_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_187_),
  .S(_188_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_170_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_169_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_168_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_167_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_166_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_165_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_164_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_163_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_162_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_161_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$4dc5718e86f31fe555f7d39cf5ab7078c09f577a\dctu

module \$paramod$53ab2e60687d01e7461fdffe1d34a14bacda6928\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _057_ (
  .A(y[0]),
  .ZN(_047_)
);

INV_X1 _058_ (
  .A(y[1]),
  .ZN(_048_)
);

INV_X1 _059_ (
  .A(_051_),
  .ZN(_008_)
);

BUF_X4 _060_ (
  .A(y[2]),
  .Z(_009_)
);

NAND2_X1 _061_ (
  .A1(_008_),
  .A2(_009_),
  .ZN(_010_)
);

INV_X4 _062_ (
  .A(_009_),
  .ZN(_011_)
);

NAND2_X1 _063_ (
  .A1(_011_),
  .A2(_053_),
  .ZN(_012_)
);

BUF_X4 _064_ (
  .A(ena),
  .Z(_013_)
);

NAND3_X1 _065_ (
  .A1(_010_),
  .A2(_012_),
  .A3(_013_),
  .ZN(_014_)
);

INV_X4 _066_ (
  .A(_013_),
  .ZN(_015_)
);

BUF_X16 _067_ (
  .A(_015_),
  .Z(_016_)
);

NAND2_X1 _068_ (
  .A1(_016_),
  .A2(\coef[13] ),
  .ZN(_017_)
);

NAND2_X1 _069_ (
  .A1(_014_),
  .A2(_017_),
  .ZN(_000_)
);

INV_X1 _070_ (
  .A(_050_),
  .ZN(_018_)
);

NAND2_X1 _071_ (
  .A1(_011_),
  .A2(_018_),
  .ZN(_019_)
);

NAND2_X1 _072_ (
  .A1(_009_),
  .A2(_050_),
  .ZN(_020_)
);

NAND3_X1 _073_ (
  .A1(_019_),
  .A2(_013_),
  .A3(_020_),
  .ZN(_021_)
);

NAND2_X1 _074_ (
  .A1(_016_),
  .A2(\coef[14] ),
  .ZN(_022_)
);

NAND2_X1 _075_ (
  .A1(_021_),
  .A2(_022_),
  .ZN(_001_)
);

NAND2_X2 _076_ (
  .A1(_016_),
  .A2(\coef[15] ),
  .ZN(_023_)
);

OAI21_X2 _077_ (
  .A(_023_),
  .B1(y[1]),
  .B2(_016_),
  .ZN(_002_)
);

NAND2_X2 _078_ (
  .A1(_016_),
  .A2(\coef[12] ),
  .ZN(_024_)
);

OAI21_X2 _079_ (
  .A(_024_),
  .B1(_011_),
  .B2(_016_),
  .ZN(_003_)
);

INV_X1 _080_ (
  .A(_049_),
  .ZN(_025_)
);

NAND2_X1 _081_ (
  .A1(_025_),
  .A2(_009_),
  .ZN(_026_)
);

NAND2_X1 _082_ (
  .A1(_011_),
  .A2(_055_),
  .ZN(_027_)
);

NAND3_X1 _083_ (
  .A1(_026_),
  .A2(_027_),
  .A3(_013_),
  .ZN(_028_)
);

NAND2_X1 _084_ (
  .A1(_016_),
  .A2(\coef[21] ),
  .ZN(_029_)
);

NAND2_X1 _085_ (
  .A1(_028_),
  .A2(_029_),
  .ZN(_004_)
);

NAND2_X1 _086_ (
  .A1(_018_),
  .A2(_009_),
  .ZN(_030_)
);

NAND2_X1 _087_ (
  .A1(_011_),
  .A2(_050_),
  .ZN(_031_)
);

NAND3_X1 _088_ (
  .A1(_030_),
  .A2(_031_),
  .A3(_013_),
  .ZN(_032_)
);

NAND2_X1 _089_ (
  .A1(_016_),
  .A2(\coef[22] ),
  .ZN(_033_)
);

NAND2_X1 _090_ (
  .A1(_032_),
  .A2(_033_),
  .ZN(_005_)
);

NAND2_X2 _091_ (
  .A1(_016_),
  .A2(\coef[23] ),
  .ZN(_034_)
);

OAI21_X2 _092_ (
  .A(_034_),
  .B1(_047_),
  .B2(_016_),
  .ZN(_006_)
);

NAND2_X1 _093_ (
  .A1(_015_),
  .A2(\coef[28] ),
  .ZN(_035_)
);

NAND2_X1 _094_ (
  .A1(_009_),
  .A2(_053_),
  .ZN(_036_)
);

NAND2_X1 _095_ (
  .A1(_036_),
  .A2(_013_),
  .ZN(_037_)
);

NOR2_X1 _096_ (
  .A1(_009_),
  .A2(_051_),
  .ZN(_038_)
);

OAI21_X1 _097_ (
  .A(_035_),
  .B1(_037_),
  .B2(_038_),
  .ZN(_007_)
);

HA_X1 _098_ (
  .A(_047_),
  .B(_048_),
  .CO(_049_),
  .S(_050_)
);

HA_X1 _099_ (
  .A(_047_),
  .B(y[1]),
  .CO(_051_),
  .S(_052_)
);

HA_X1 _100_ (
  .A(y[0]),
  .B(_048_),
  .CO(_053_),
  .S(_054_)
);

HA_X1 _101_ (
  .A(y[0]),
  .B(y[1]),
  .CO(_055_),
  .S(_056_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_042_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_041_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_040_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_045_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_046_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_039_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_044_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_043_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$53ab2e60687d01e7461fdffe1d34a14bacda6928\dctu

module \$paramod$56b31b71c3bccc1fb1f134779b3bdd5ab1b461c7\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _193_ (
  .A(x[0]),
  .ZN(_175_)
);

INV_X1 _194_ (
  .A(x[1]),
  .ZN(_176_)
);

INV_X2 _195_ (
  .A(x[2]),
  .ZN(_106_)
);

BUF_X8 _196_ (
  .A(_106_),
  .Z(_107_)
);

NAND2_X4 _197_ (
  .A1(_107_),
  .A2(_177_),
  .ZN(_108_)
);

INV_X1 _198_ (
  .A(_191_),
  .ZN(_109_)
);

BUF_X4 _199_ (
  .A(x[2]),
  .Z(_110_)
);

NAND2_X2 _200_ (
  .A1(_109_),
  .A2(_110_),
  .ZN(_111_)
);

BUF_X4 _201_ (
  .A(y[0]),
  .Z(_112_)
);

BUF_X4 _202_ (
  .A(_112_),
  .Z(_113_)
);

NAND3_X1 _203_ (
  .A1(_108_),
  .A2(_111_),
  .A3(_113_),
  .ZN(_114_)
);

NAND2_X1 _204_ (
  .A1(_106_),
  .A2(_178_),
  .ZN(_115_)
);

INV_X1 _205_ (
  .A(_178_),
  .ZN(_116_)
);

NAND2_X1 _206_ (
  .A1(_116_),
  .A2(x[2]),
  .ZN(_117_)
);

INV_X8 _207_ (
  .A(_112_),
  .ZN(_118_)
);

BUF_X8 _208_ (
  .A(_118_),
  .Z(_119_)
);

NAND3_X1 _209_ (
  .A1(_115_),
  .A2(_117_),
  .A3(_119_),
  .ZN(_120_)
);

NAND2_X1 _210_ (
  .A1(_114_),
  .A2(_120_),
  .ZN(_121_)
);

BUF_X4 _211_ (
  .A(y[1]),
  .Z(_122_)
);

INV_X2 _212_ (
  .A(_122_),
  .ZN(_123_)
);

BUF_X2 _213_ (
  .A(_123_),
  .Z(_124_)
);

NAND2_X1 _214_ (
  .A1(_121_),
  .A2(_124_),
  .ZN(_125_)
);

INV_X1 _215_ (
  .A(_187_),
  .ZN(_126_)
);

NAND2_X2 _216_ (
  .A1(_107_),
  .A2(_126_),
  .ZN(_127_)
);

NAND2_X2 _217_ (
  .A1(_110_),
  .A2(_181_),
  .ZN(_128_)
);

NAND3_X2 _218_ (
  .A1(_127_),
  .A2(_119_),
  .A3(_128_),
  .ZN(_129_)
);

NAND2_X1 _219_ (
  .A1(_176_),
  .A2(_113_),
  .ZN(_130_)
);

NAND2_X1 _220_ (
  .A1(_129_),
  .A2(_130_),
  .ZN(_131_)
);

BUF_X2 _221_ (
  .A(_122_),
  .Z(_132_)
);

NAND2_X1 _222_ (
  .A1(_131_),
  .A2(_132_),
  .ZN(_133_)
);

BUF_X2 _223_ (
  .A(y[2]),
  .Z(_134_)
);

INV_X1 _224_ (
  .A(_134_),
  .ZN(_135_)
);

NAND3_X1 _225_ (
  .A1(_125_),
  .A2(_133_),
  .A3(_135_),
  .ZN(_136_)
);

NAND2_X2 _226_ (
  .A1(_107_),
  .A2(_185_),
  .ZN(_137_)
);

INV_X1 _227_ (
  .A(_183_),
  .ZN(_138_)
);

NAND2_X2 _228_ (
  .A1(_138_),
  .A2(_110_),
  .ZN(_139_)
);

NAND2_X1 _229_ (
  .A1(_137_),
  .A2(_139_),
  .ZN(_140_)
);

NAND2_X1 _230_ (
  .A1(_140_),
  .A2(_113_),
  .ZN(_141_)
);

AOI21_X2 _231_ (
  .A(_122_),
  .B1(_119_),
  .B2(_176_),
  .ZN(_142_)
);

AOI21_X1 _232_ (
  .A(_135_),
  .B1(_141_),
  .B2(_142_),
  .ZN(_143_)
);

INV_X1 _233_ (
  .A(_179_),
  .ZN(_144_)
);

NAND2_X4 _234_ (
  .A1(_107_),
  .A2(_144_),
  .ZN(_145_)
);

NAND2_X4 _235_ (
  .A1(_110_),
  .A2(_189_),
  .ZN(_146_)
);

NAND2_X1 _236_ (
  .A1(_145_),
  .A2(_146_),
  .ZN(_147_)
);

NAND2_X1 _237_ (
  .A1(_147_),
  .A2(_119_),
  .ZN(_148_)
);

NAND3_X2 _238_ (
  .A1(_115_),
  .A2(_117_),
  .A3(_112_),
  .ZN(_149_)
);

NAND3_X1 _239_ (
  .A1(_148_),
  .A2(_149_),
  .A3(_132_),
  .ZN(_150_)
);

NAND2_X1 _240_ (
  .A1(_143_),
  .A2(_150_),
  .ZN(_151_)
);

BUF_X2 _241_ (
  .A(ena),
  .Z(_152_)
);

NAND3_X1 _242_ (
  .A1(_136_),
  .A2(_151_),
  .A3(_152_),
  .ZN(_153_)
);

INV_X1 _243_ (
  .A(_152_),
  .ZN(_154_)
);

NAND2_X1 _244_ (
  .A1(_154_),
  .A2(\coef[21] ),
  .ZN(_155_)
);

NAND2_X1 _245_ (
  .A1(_153_),
  .A2(_155_),
  .ZN(_000_)
);

NAND3_X1 _246_ (
  .A1(_137_),
  .A2(_139_),
  .A3(_119_),
  .ZN(_156_)
);

NAND3_X1 _247_ (
  .A1(_114_),
  .A2(_156_),
  .A3(_132_),
  .ZN(_157_)
);

NAND2_X2 _248_ (
  .A1(_107_),
  .A2(_116_),
  .ZN(_158_)
);

NAND2_X4 _249_ (
  .A1(_110_),
  .A2(_178_),
  .ZN(_159_)
);

NAND3_X4 _250_ (
  .A1(_158_),
  .A2(_118_),
  .A3(_159_),
  .ZN(_160_)
);

NAND3_X1 _251_ (
  .A1(_149_),
  .A2(_160_),
  .A3(_123_),
  .ZN(_161_)
);

NAND3_X1 _252_ (
  .A1(_157_),
  .A2(_161_),
  .A3(_135_),
  .ZN(_162_)
);

NAND3_X1 _253_ (
  .A1(_145_),
  .A2(_119_),
  .A3(_146_),
  .ZN(_163_)
);

NAND3_X1 _254_ (
  .A1(_127_),
  .A2(_113_),
  .A3(_128_),
  .ZN(_164_)
);

NAND3_X1 _255_ (
  .A1(_163_),
  .A2(_164_),
  .A3(_123_),
  .ZN(_165_)
);

NAND3_X1 _256_ (
  .A1(_149_),
  .A2(_160_),
  .A3(_122_),
  .ZN(_009_)
);

NAND3_X1 _257_ (
  .A1(_165_),
  .A2(_009_),
  .A3(_134_),
  .ZN(_010_)
);

NAND2_X1 _258_ (
  .A1(_162_),
  .A2(_010_),
  .ZN(_011_)
);

NAND2_X1 _259_ (
  .A1(_011_),
  .A2(_152_),
  .ZN(_012_)
);

NAND2_X1 _260_ (
  .A1(_154_),
  .A2(\coef[23] ),
  .ZN(_013_)
);

NAND2_X1 _261_ (
  .A1(_012_),
  .A2(_013_),
  .ZN(_001_)
);

NAND3_X2 _262_ (
  .A1(_108_),
  .A2(_111_),
  .A3(_118_),
  .ZN(_014_)
);

NAND3_X1 _263_ (
  .A1(_149_),
  .A2(_014_),
  .A3(_132_),
  .ZN(_015_)
);

NAND2_X1 _264_ (
  .A1(_144_),
  .A2(_110_),
  .ZN(_016_)
);

NAND2_X1 _265_ (
  .A1(_107_),
  .A2(_189_),
  .ZN(_017_)
);

NAND3_X2 _266_ (
  .A1(_016_),
  .A2(_017_),
  .A3(_118_),
  .ZN(_018_)
);

NAND2_X1 _267_ (
  .A1(x[0]),
  .A2(_112_),
  .ZN(_019_)
);

NAND3_X1 _268_ (
  .A1(_018_),
  .A2(_123_),
  .A3(_019_),
  .ZN(_020_)
);

NAND3_X1 _269_ (
  .A1(_015_),
  .A2(_020_),
  .A3(_134_),
  .ZN(_021_)
);

NAND3_X2 _270_ (
  .A1(_145_),
  .A2(_112_),
  .A3(_146_),
  .ZN(_022_)
);

NAND3_X1 _271_ (
  .A1(_160_),
  .A2(_022_),
  .A3(_123_),
  .ZN(_023_)
);

NAND2_X1 _272_ (
  .A1(_107_),
  .A2(_109_),
  .ZN(_024_)
);

NAND2_X1 _273_ (
  .A1(_110_),
  .A2(_177_),
  .ZN(_025_)
);

NAND3_X2 _274_ (
  .A1(_024_),
  .A2(_113_),
  .A3(_025_),
  .ZN(_026_)
);

NOR2_X1 _275_ (
  .A1(x[0]),
  .A2(_112_),
  .ZN(_027_)
);

INV_X1 _276_ (
  .A(_027_),
  .ZN(_028_)
);

NAND3_X1 _277_ (
  .A1(_026_),
  .A2(_122_),
  .A3(_028_),
  .ZN(_029_)
);

NAND3_X1 _278_ (
  .A1(_023_),
  .A2(_029_),
  .A3(_135_),
  .ZN(_030_)
);

NAND2_X1 _279_ (
  .A1(_021_),
  .A2(_030_),
  .ZN(_031_)
);

NAND2_X1 _280_ (
  .A1(_031_),
  .A2(_152_),
  .ZN(_032_)
);

NAND2_X1 _281_ (
  .A1(_154_),
  .A2(\coef[24] ),
  .ZN(_033_)
);

NAND2_X1 _282_ (
  .A1(_032_),
  .A2(_033_),
  .ZN(_002_)
);

NOR2_X1 _283_ (
  .A1(_112_),
  .A2(_110_),
  .ZN(_034_)
);

INV_X1 _284_ (
  .A(_034_),
  .ZN(_035_)
);

NAND2_X1 _285_ (
  .A1(_149_),
  .A2(_035_),
  .ZN(_036_)
);

NAND2_X1 _286_ (
  .A1(_036_),
  .A2(_124_),
  .ZN(_037_)
);

NAND3_X1 _287_ (
  .A1(_028_),
  .A2(_122_),
  .A3(_130_),
  .ZN(_038_)
);

NAND3_X1 _288_ (
  .A1(_037_),
  .A2(_134_),
  .A3(_038_),
  .ZN(_039_)
);

OAI21_X1 _289_ (
  .A(_019_),
  .B1(_176_),
  .B2(_113_),
  .ZN(_040_)
);

NAND2_X1 _290_ (
  .A1(_040_),
  .A2(_123_),
  .ZN(_041_)
);

INV_X1 _291_ (
  .A(_160_),
  .ZN(_042_)
);

OAI21_X2 _292_ (
  .A(_122_),
  .B1(_119_),
  .B2(_107_),
  .ZN(_043_)
);

OAI21_X1 _293_ (
  .A(_041_),
  .B1(_042_),
  .B2(_043_),
  .ZN(_044_)
);

NAND2_X1 _294_ (
  .A1(_044_),
  .A2(_135_),
  .ZN(_045_)
);

NAND2_X1 _295_ (
  .A1(_039_),
  .A2(_045_),
  .ZN(_046_)
);

NAND2_X1 _296_ (
  .A1(_046_),
  .A2(_152_),
  .ZN(_047_)
);

NAND2_X1 _297_ (
  .A1(_154_),
  .A2(\coef[10] ),
  .ZN(_048_)
);

NAND2_X1 _298_ (
  .A1(_047_),
  .A2(_048_),
  .ZN(_003_)
);

NAND2_X1 _299_ (
  .A1(_149_),
  .A2(_156_),
  .ZN(_049_)
);

NAND2_X1 _300_ (
  .A1(_049_),
  .A2(_124_),
  .ZN(_050_)
);

NAND2_X1 _301_ (
  .A1(x[1]),
  .A2(_113_),
  .ZN(_051_)
);

NAND2_X1 _302_ (
  .A1(_129_),
  .A2(_051_),
  .ZN(_052_)
);

NAND2_X1 _303_ (
  .A1(_052_),
  .A2(_132_),
  .ZN(_053_)
);

NAND3_X1 _304_ (
  .A1(_050_),
  .A2(_053_),
  .A3(_134_),
  .ZN(_054_)
);

NAND3_X1 _305_ (
  .A1(_160_),
  .A2(_164_),
  .A3(_122_),
  .ZN(_055_)
);

NAND3_X1 _306_ (
  .A1(_137_),
  .A2(_139_),
  .A3(_113_),
  .ZN(_056_)
);

NAND2_X1 _307_ (
  .A1(_056_),
  .A2(_142_),
  .ZN(_057_)
);

NAND2_X1 _308_ (
  .A1(_055_),
  .A2(_057_),
  .ZN(_058_)
);

NAND2_X1 _309_ (
  .A1(_058_),
  .A2(_135_),
  .ZN(_059_)
);

NAND3_X1 _310_ (
  .A1(_054_),
  .A2(_059_),
  .A3(_152_),
  .ZN(_060_)
);

NAND2_X1 _311_ (
  .A1(_154_),
  .A2(\coef[26] ),
  .ZN(_061_)
);

NAND2_X1 _312_ (
  .A1(_060_),
  .A2(_061_),
  .ZN(_004_)
);

NOR2_X1 _313_ (
  .A1(_152_),
  .A2(\coef[13] ),
  .ZN(_062_)
);

INV_X1 _314_ (
  .A(_043_),
  .ZN(_063_)
);

AOI21_X1 _315_ (
  .A(_134_),
  .B1(_018_),
  .B2(_063_),
  .ZN(_064_)
);

NAND2_X2 _316_ (
  .A1(_107_),
  .A2(_138_),
  .ZN(_065_)
);

NAND2_X1 _317_ (
  .A1(_110_),
  .A2(_185_),
  .ZN(_066_)
);

NAND3_X1 _318_ (
  .A1(_065_),
  .A2(_113_),
  .A3(_066_),
  .ZN(_067_)
);

NAND3_X1 _319_ (
  .A1(_067_),
  .A2(_124_),
  .A3(_028_),
  .ZN(_068_)
);

AOI21_X1 _320_ (
  .A(_154_),
  .B1(_064_),
  .B2(_068_),
  .ZN(_069_)
);

NAND2_X1 _321_ (
  .A1(_107_),
  .A2(_181_),
  .ZN(_070_)
);

NAND2_X1 _322_ (
  .A1(_126_),
  .A2(_110_),
  .ZN(_071_)
);

NAND3_X1 _323_ (
  .A1(_070_),
  .A2(_071_),
  .A3(_119_),
  .ZN(_072_)
);

NAND3_X1 _324_ (
  .A1(_072_),
  .A2(_132_),
  .A3(_019_),
  .ZN(_073_)
);

NAND3_X1 _325_ (
  .A1(_026_),
  .A2(_124_),
  .A3(_035_),
  .ZN(_074_)
);

NAND3_X1 _326_ (
  .A1(_073_),
  .A2(_074_),
  .A3(_134_),
  .ZN(_075_)
);

AOI21_X2 _327_ (
  .A(_062_),
  .B1(_069_),
  .B2(_075_),
  .ZN(_005_)
);

NAND3_X1 _328_ (
  .A1(_056_),
  .A2(_014_),
  .A3(_132_),
  .ZN(_076_)
);

NAND3_X1 _329_ (
  .A1(_070_),
  .A2(_071_),
  .A3(_113_),
  .ZN(_077_)
);

NAND3_X1 _330_ (
  .A1(_018_),
  .A2(_077_),
  .A3(_123_),
  .ZN(_078_)
);

NAND3_X1 _331_ (
  .A1(_076_),
  .A2(_078_),
  .A3(_134_),
  .ZN(_079_)
);

NAND3_X1 _332_ (
  .A1(_129_),
  .A2(_022_),
  .A3(_123_),
  .ZN(_080_)
);

NAND3_X1 _333_ (
  .A1(_065_),
  .A2(_119_),
  .A3(_066_),
  .ZN(_081_)
);

NAND3_X1 _334_ (
  .A1(_026_),
  .A2(_081_),
  .A3(_122_),
  .ZN(_082_)
);

NAND3_X1 _335_ (
  .A1(_080_),
  .A2(_082_),
  .A3(_135_),
  .ZN(_083_)
);

NAND2_X1 _336_ (
  .A1(_079_),
  .A2(_083_),
  .ZN(_084_)
);

NAND2_X1 _337_ (
  .A1(_084_),
  .A2(_152_),
  .ZN(_085_)
);

NAND2_X1 _338_ (
  .A1(_154_),
  .A2(\coef[28] ),
  .ZN(_086_)
);

NAND2_X1 _339_ (
  .A1(_085_),
  .A2(_086_),
  .ZN(_006_)
);

NAND2_X1 _340_ (
  .A1(_072_),
  .A2(_022_),
  .ZN(_087_)
);

NAND2_X1 _341_ (
  .A1(_087_),
  .A2(_124_),
  .ZN(_088_)
);

NAND2_X1 _342_ (
  .A1(_176_),
  .A2(_119_),
  .ZN(_089_)
);

NAND3_X1 _343_ (
  .A1(_089_),
  .A2(_132_),
  .A3(_019_),
  .ZN(_090_)
);

NAND3_X1 _344_ (
  .A1(_088_),
  .A2(_135_),
  .A3(_090_),
  .ZN(_091_)
);

NAND2_X1 _345_ (
  .A1(_014_),
  .A2(_067_),
  .ZN(_092_)
);

NAND2_X1 _346_ (
  .A1(_092_),
  .A2(_132_),
  .ZN(_093_)
);

NAND3_X1 _347_ (
  .A1(_028_),
  .A2(_124_),
  .A3(_051_),
  .ZN(_094_)
);

NAND3_X1 _348_ (
  .A1(_093_),
  .A2(_134_),
  .A3(_094_),
  .ZN(_095_)
);

NAND3_X1 _349_ (
  .A1(_091_),
  .A2(_095_),
  .A3(_152_),
  .ZN(_096_)
);

NAND2_X1 _350_ (
  .A1(_154_),
  .A2(\coef[29] ),
  .ZN(_097_)
);

NAND2_X1 _351_ (
  .A1(_096_),
  .A2(_097_),
  .ZN(_007_)
);

NOR2_X1 _352_ (
  .A1(_152_),
  .A2(\coef[30] ),
  .ZN(_098_)
);

NAND3_X1 _353_ (
  .A1(_014_),
  .A2(_022_),
  .A3(_124_),
  .ZN(_099_)
);

AOI21_X1 _354_ (
  .A(_134_),
  .B1(_147_),
  .B2(_132_),
  .ZN(_100_)
);

AOI21_X1 _355_ (
  .A(_154_),
  .B1(_099_),
  .B2(_100_),
  .ZN(_101_)
);

NAND2_X1 _356_ (
  .A1(_108_),
  .A2(_111_),
  .ZN(_102_)
);

AOI21_X1 _357_ (
  .A(_135_),
  .B1(_102_),
  .B2(_124_),
  .ZN(_103_)
);

NAND2_X1 _358_ (
  .A1(_014_),
  .A2(_022_),
  .ZN(_104_)
);

OAI21_X1 _359_ (
  .A(_103_),
  .B1(_104_),
  .B2(_124_),
  .ZN(_105_)
);

AOI21_X1 _360_ (
  .A(_098_),
  .B1(_101_),
  .B2(_105_),
  .ZN(_008_)
);

HA_X1 _361_ (
  .A(_175_),
  .B(_176_),
  .CO(_177_),
  .S(_178_)
);

HA_X1 _362_ (
  .A(_175_),
  .B(_176_),
  .CO(_179_),
  .S(_180_)
);

HA_X1 _363_ (
  .A(_175_),
  .B(x[1]),
  .CO(_181_),
  .S(_182_)
);

HA_X1 _364_ (
  .A(_175_),
  .B(x[1]),
  .CO(_183_),
  .S(_184_)
);

HA_X1 _365_ (
  .A(x[0]),
  .B(_176_),
  .CO(_185_),
  .S(_186_)
);

HA_X1 _366_ (
  .A(x[0]),
  .B(_176_),
  .CO(_187_),
  .S(_188_)
);

HA_X1 _367_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_189_),
  .S(_190_)
);

HA_X1 _368_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_191_),
  .S(_192_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_174_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_173_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_172_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_171_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_170_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_169_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_168_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_167_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_166_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$56b31b71c3bccc1fb1f134779b3bdd5ab1b461c7\dctu

module \$paramod$5778094f610ca183dd46956f589e4ea513d2316c\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _181_ (
  .A(x[1]),
  .ZN(_164_)
);

INV_X1 _182_ (
  .A(x[0]),
  .ZN(_163_)
);

BUF_X2 _183_ (
  .A(y[2]),
  .Z(_094_)
);

INV_X2 _184_ (
  .A(_094_),
  .ZN(_095_)
);

BUF_X2 _185_ (
  .A(y[1]),
  .Z(_096_)
);

BUF_X2 _186_ (
  .A(_096_),
  .Z(_097_)
);

BUF_X4 _187_ (
  .A(x[2]),
  .Z(_098_)
);

XNOR2_X2 _188_ (
  .A(_098_),
  .B(_166_),
  .ZN(_099_)
);

INV_X2 _189_ (
  .A(_099_),
  .ZN(_100_)
);

BUF_X4 _190_ (
  .A(y[0]),
  .Z(_101_)
);

BUF_X4 _191_ (
  .A(_101_),
  .Z(_102_)
);

NAND2_X4 _192_ (
  .A1(_100_),
  .A2(_102_),
  .ZN(_103_)
);

INV_X4 _193_ (
  .A(_098_),
  .ZN(_104_)
);

NAND2_X2 _194_ (
  .A1(_104_),
  .A2(_173_),
  .ZN(_105_)
);

INV_X1 _195_ (
  .A(_171_),
  .ZN(_106_)
);

BUF_X16 _196_ (
  .A(_098_),
  .Z(_107_)
);

NAND2_X4 _197_ (
  .A1(_106_),
  .A2(_107_),
  .ZN(_108_)
);

NAND2_X2 _198_ (
  .A1(_105_),
  .A2(_108_),
  .ZN(_109_)
);

INV_X8 _199_ (
  .A(_101_),
  .ZN(_110_)
);

BUF_X8 _200_ (
  .A(_110_),
  .Z(_111_)
);

NAND2_X1 _201_ (
  .A1(_109_),
  .A2(_111_),
  .ZN(_112_)
);

AOI21_X2 _202_ (
  .A(_097_),
  .B1(_103_),
  .B2(_112_),
  .ZN(_113_)
);

INV_X1 _203_ (
  .A(_167_),
  .ZN(_114_)
);

NAND2_X2 _204_ (
  .A1(_104_),
  .A2(_114_),
  .ZN(_115_)
);

NAND2_X4 _205_ (
  .A1(_107_),
  .A2(_177_),
  .ZN(_116_)
);

NAND3_X1 _206_ (
  .A1(_115_),
  .A2(_102_),
  .A3(_116_),
  .ZN(_117_)
);

NAND2_X2 _207_ (
  .A1(_110_),
  .A2(x[1]),
  .ZN(_118_)
);

NAND3_X1 _208_ (
  .A1(_117_),
  .A2(_097_),
  .A3(_118_),
  .ZN(_119_)
);

INV_X1 _209_ (
  .A(_119_),
  .ZN(_120_)
);

OAI21_X1 _210_ (
  .A(_095_),
  .B1(_113_),
  .B2(_120_),
  .ZN(_121_)
);

BUF_X2 _211_ (
  .A(ena),
  .Z(_122_)
);

INV_X1 _212_ (
  .A(_122_),
  .ZN(_123_)
);

NAND2_X2 _213_ (
  .A1(_099_),
  .A2(_110_),
  .ZN(_124_)
);

INV_X1 _214_ (
  .A(_175_),
  .ZN(_125_)
);

NAND2_X2 _215_ (
  .A1(_104_),
  .A2(_125_),
  .ZN(_126_)
);

NAND2_X1 _216_ (
  .A1(_098_),
  .A2(_169_),
  .ZN(_127_)
);

NAND2_X1 _217_ (
  .A1(_126_),
  .A2(_127_),
  .ZN(_128_)
);

NAND2_X1 _218_ (
  .A1(_128_),
  .A2(_102_),
  .ZN(_129_)
);

NAND3_X1 _219_ (
  .A1(_124_),
  .A2(_129_),
  .A3(_097_),
  .ZN(_130_)
);

NAND2_X2 _220_ (
  .A1(_104_),
  .A2(_165_),
  .ZN(_131_)
);

INV_X1 _221_ (
  .A(_179_),
  .ZN(_132_)
);

NAND2_X4 _222_ (
  .A1(_132_),
  .A2(_107_),
  .ZN(_133_)
);

NAND3_X1 _223_ (
  .A1(_131_),
  .A2(_133_),
  .A3(_111_),
  .ZN(_134_)
);

NAND2_X1 _224_ (
  .A1(_164_),
  .A2(_101_),
  .ZN(_135_)
);

NAND2_X1 _225_ (
  .A1(_135_),
  .A2(_094_),
  .ZN(_136_)
);

INV_X1 _226_ (
  .A(_136_),
  .ZN(_137_)
);

NAND2_X1 _227_ (
  .A1(_134_),
  .A2(_137_),
  .ZN(_138_)
);

NAND2_X1 _228_ (
  .A1(_096_),
  .A2(_094_),
  .ZN(_139_)
);

NAND2_X1 _229_ (
  .A1(_138_),
  .A2(_139_),
  .ZN(_140_)
);

AOI21_X1 _230_ (
  .A(_123_),
  .B1(_130_),
  .B2(_140_),
  .ZN(_141_)
);

NAND2_X1 _231_ (
  .A1(_121_),
  .A2(_141_),
  .ZN(_142_)
);

NAND2_X1 _232_ (
  .A1(_123_),
  .A2(\coef[21] ),
  .ZN(_143_)
);

NAND2_X1 _233_ (
  .A1(_142_),
  .A2(_143_),
  .ZN(_000_)
);

NAND3_X2 _234_ (
  .A1(_131_),
  .A2(_133_),
  .A3(_096_),
  .ZN(_144_)
);

INV_X2 _235_ (
  .A(_096_),
  .ZN(_145_)
);

NAND3_X1 _236_ (
  .A1(_126_),
  .A2(_145_),
  .A3(_127_),
  .ZN(_146_)
);

NAND3_X1 _237_ (
  .A1(_144_),
  .A2(_146_),
  .A3(_102_),
  .ZN(_147_)
);

NAND3_X1 _238_ (
  .A1(_147_),
  .A2(_095_),
  .A3(_118_),
  .ZN(_148_)
);

NAND3_X1 _239_ (
  .A1(_115_),
  .A2(_145_),
  .A3(_116_),
  .ZN(_149_)
);

NAND2_X1 _240_ (
  .A1(_149_),
  .A2(_111_),
  .ZN(_150_)
);

NOR2_X1 _241_ (
  .A1(_109_),
  .A2(_145_),
  .ZN(_151_)
);

OAI21_X1 _242_ (
  .A(_137_),
  .B1(_150_),
  .B2(_151_),
  .ZN(_152_)
);

NAND2_X1 _243_ (
  .A1(_148_),
  .A2(_152_),
  .ZN(_153_)
);

NAND2_X1 _244_ (
  .A1(_153_),
  .A2(_122_),
  .ZN(_009_)
);

NAND2_X1 _245_ (
  .A1(_123_),
  .A2(\coef[23] ),
  .ZN(_010_)
);

NAND2_X1 _246_ (
  .A1(_009_),
  .A2(_010_),
  .ZN(_001_)
);

NAND2_X1 _247_ (
  .A1(_104_),
  .A2(_169_),
  .ZN(_011_)
);

NAND2_X2 _248_ (
  .A1(_125_),
  .A2(_107_),
  .ZN(_012_)
);

NAND3_X1 _249_ (
  .A1(_011_),
  .A2(_012_),
  .A3(_111_),
  .ZN(_013_)
);

NAND3_X4 _250_ (
  .A1(_105_),
  .A2(_108_),
  .A3(_102_),
  .ZN(_014_)
);

NAND2_X1 _251_ (
  .A1(_013_),
  .A2(_014_),
  .ZN(_015_)
);

NAND2_X1 _252_ (
  .A1(_015_),
  .A2(_097_),
  .ZN(_016_)
);

NAND2_X1 _253_ (
  .A1(_104_),
  .A2(_111_),
  .ZN(_017_)
);

NAND3_X1 _254_ (
  .A1(_017_),
  .A2(_135_),
  .A3(_145_),
  .ZN(_018_)
);

NAND3_X1 _255_ (
  .A1(_016_),
  .A2(_094_),
  .A3(_018_),
  .ZN(_019_)
);

NAND3_X2 _256_ (
  .A1(_126_),
  .A2(_110_),
  .A3(_127_),
  .ZN(_020_)
);

NAND2_X1 _257_ (
  .A1(_104_),
  .A2(_106_),
  .ZN(_021_)
);

NAND2_X2 _258_ (
  .A1(_107_),
  .A2(_173_),
  .ZN(_022_)
);

NAND3_X1 _259_ (
  .A1(_021_),
  .A2(_102_),
  .A3(_022_),
  .ZN(_023_)
);

NAND2_X1 _260_ (
  .A1(_020_),
  .A2(_023_),
  .ZN(_024_)
);

NAND2_X1 _261_ (
  .A1(_024_),
  .A2(_145_),
  .ZN(_025_)
);

NAND2_X1 _262_ (
  .A1(_107_),
  .A2(_102_),
  .ZN(_026_)
);

NAND3_X1 _263_ (
  .A1(_118_),
  .A2(_026_),
  .A3(_097_),
  .ZN(_027_)
);

NAND3_X1 _264_ (
  .A1(_025_),
  .A2(_095_),
  .A3(_027_),
  .ZN(_028_)
);

NAND3_X1 _265_ (
  .A1(_019_),
  .A2(_028_),
  .A3(_122_),
  .ZN(_029_)
);

NAND2_X1 _266_ (
  .A1(_123_),
  .A2(\coef[24] ),
  .ZN(_030_)
);

NAND2_X1 _267_ (
  .A1(_029_),
  .A2(_030_),
  .ZN(_002_)
);

NOR2_X1 _268_ (
  .A1(_122_),
  .A2(\coef[10] ),
  .ZN(_031_)
);

NAND2_X1 _269_ (
  .A1(_118_),
  .A2(_094_),
  .ZN(_032_)
);

INV_X1 _270_ (
  .A(_032_),
  .ZN(_033_)
);

NAND2_X4 _271_ (
  .A1(_103_),
  .A2(_033_),
  .ZN(_034_)
);

NAND2_X4 _272_ (
  .A1(_034_),
  .A2(_139_),
  .ZN(_035_)
);

NAND2_X1 _273_ (
  .A1(_111_),
  .A2(_163_),
  .ZN(_036_)
);

NAND3_X1 _274_ (
  .A1(_036_),
  .A2(_097_),
  .A3(_026_),
  .ZN(_037_)
);

AOI21_X2 _275_ (
  .A(_123_),
  .B1(_035_),
  .B2(_037_),
  .ZN(_038_)
);

NAND2_X1 _276_ (
  .A1(_124_),
  .A2(_135_),
  .ZN(_039_)
);

NAND2_X1 _277_ (
  .A1(_039_),
  .A2(_097_),
  .ZN(_040_)
);

NAND2_X2 _278_ (
  .A1(_110_),
  .A2(_107_),
  .ZN(_041_)
);

NAND2_X1 _279_ (
  .A1(_163_),
  .A2(_102_),
  .ZN(_042_)
);

NAND2_X1 _280_ (
  .A1(_041_),
  .A2(_042_),
  .ZN(_043_)
);

NAND2_X1 _281_ (
  .A1(_043_),
  .A2(_145_),
  .ZN(_044_)
);

NAND3_X1 _282_ (
  .A1(_040_),
  .A2(_095_),
  .A3(_044_),
  .ZN(_045_)
);

AOI21_X2 _283_ (
  .A(_031_),
  .B1(_038_),
  .B2(_045_),
  .ZN(_003_)
);

AOI21_X4 _284_ (
  .A(_123_),
  .B1(_035_),
  .B2(_144_),
  .ZN(_046_)
);

NAND3_X1 _285_ (
  .A1(_040_),
  .A2(_095_),
  .A3(_149_),
  .ZN(_047_)
);

NAND2_X2 _286_ (
  .A1(_046_),
  .A2(_047_),
  .ZN(_048_)
);

NAND2_X1 _287_ (
  .A1(_123_),
  .A2(\coef[26] ),
  .ZN(_049_)
);

NAND2_X2 _288_ (
  .A1(_048_),
  .A2(_049_),
  .ZN(_004_)
);

NOR2_X1 _289_ (
  .A1(_122_),
  .A2(\coef[13] ),
  .ZN(_050_)
);

NAND2_X1 _290_ (
  .A1(_104_),
  .A2(_179_),
  .ZN(_051_)
);

INV_X1 _291_ (
  .A(_165_),
  .ZN(_052_)
);

NAND2_X2 _292_ (
  .A1(_052_),
  .A2(_107_),
  .ZN(_053_)
);

NAND2_X4 _293_ (
  .A1(_051_),
  .A2(_053_),
  .ZN(_054_)
);

NAND2_X4 _294_ (
  .A1(_054_),
  .A2(_110_),
  .ZN(_055_)
);

AOI21_X1 _295_ (
  .A(_097_),
  .B1(_055_),
  .B2(_042_),
  .ZN(_056_)
);

NAND2_X1 _296_ (
  .A1(_041_),
  .A2(_096_),
  .ZN(_057_)
);

INV_X1 _297_ (
  .A(_057_),
  .ZN(_058_)
);

AND2_X2 _298_ (
  .A1(_011_),
  .A2(_012_),
  .ZN(_059_)
);

OAI21_X2 _299_ (
  .A(_058_),
  .B1(_059_),
  .B2(_111_),
  .ZN(_060_)
);

INV_X1 _300_ (
  .A(_060_),
  .ZN(_061_)
);

OAI21_X2 _301_ (
  .A(_095_),
  .B1(_056_),
  .B2(_061_),
  .ZN(_062_)
);

NOR2_X2 _302_ (
  .A1(_110_),
  .A2(_107_),
  .ZN(_063_)
);

NOR3_X1 _303_ (
  .A1(_063_),
  .A2(_096_),
  .A3(_095_),
  .ZN(_064_)
);

NAND2_X1 _304_ (
  .A1(_021_),
  .A2(_022_),
  .ZN(_065_)
);

NAND2_X1 _305_ (
  .A1(_065_),
  .A2(_111_),
  .ZN(_066_)
);

NAND2_X1 _306_ (
  .A1(_064_),
  .A2(_066_),
  .ZN(_067_)
);

NAND2_X1 _307_ (
  .A1(_067_),
  .A2(_122_),
  .ZN(_068_)
);

NAND2_X1 _308_ (
  .A1(_104_),
  .A2(_177_),
  .ZN(_069_)
);

NAND2_X2 _309_ (
  .A1(_114_),
  .A2(_107_),
  .ZN(_070_)
);

NAND3_X2 _310_ (
  .A1(_069_),
  .A2(_070_),
  .A3(_102_),
  .ZN(_071_)
);

NAND2_X1 _311_ (
  .A1(_111_),
  .A2(x[0]),
  .ZN(_072_)
);

AOI21_X1 _312_ (
  .A(_139_),
  .B1(_071_),
  .B2(_072_),
  .ZN(_073_)
);

NOR2_X1 _313_ (
  .A1(_068_),
  .A2(_073_),
  .ZN(_074_)
);

AOI21_X2 _314_ (
  .A(_050_),
  .B1(_062_),
  .B2(_074_),
  .ZN(_005_)
);

NAND3_X1 _315_ (
  .A1(_131_),
  .A2(_133_),
  .A3(_102_),
  .ZN(_075_)
);

NAND2_X2 _316_ (
  .A1(_055_),
  .A2(_075_),
  .ZN(_076_)
);

NAND2_X1 _317_ (
  .A1(_076_),
  .A2(_145_),
  .ZN(_077_)
);

NAND3_X1 _318_ (
  .A1(_016_),
  .A2(_077_),
  .A3(_094_),
  .ZN(_078_)
);

NAND3_X1 _319_ (
  .A1(_115_),
  .A2(_111_),
  .A3(_116_),
  .ZN(_079_)
);

NAND2_X1 _320_ (
  .A1(_071_),
  .A2(_079_),
  .ZN(_080_)
);

NAND2_X1 _321_ (
  .A1(_080_),
  .A2(_097_),
  .ZN(_081_)
);

NAND3_X1 _322_ (
  .A1(_025_),
  .A2(_081_),
  .A3(_095_),
  .ZN(_082_)
);

NAND3_X1 _323_ (
  .A1(_078_),
  .A2(_082_),
  .A3(_122_),
  .ZN(_083_)
);

NAND2_X1 _324_ (
  .A1(_123_),
  .A2(\coef[28] ),
  .ZN(_084_)
);

NAND2_X1 _325_ (
  .A1(_083_),
  .A2(_084_),
  .ZN(_006_)
);

NOR2_X1 _326_ (
  .A1(_122_),
  .A2(\coef[29] ),
  .ZN(_085_)
);

NAND3_X1 _327_ (
  .A1(_103_),
  .A2(_097_),
  .A3(_055_),
  .ZN(_086_)
);

NOR2_X1 _328_ (
  .A1(_063_),
  .A2(_096_),
  .ZN(_087_)
);

AOI21_X1 _329_ (
  .A(_094_),
  .B1(_020_),
  .B2(_087_),
  .ZN(_088_)
);

AOI21_X1 _330_ (
  .A(_123_),
  .B1(_086_),
  .B2(_088_),
  .ZN(_089_)
);

NAND3_X1 _331_ (
  .A1(_124_),
  .A2(_145_),
  .A3(_071_),
  .ZN(_090_)
);

AOI21_X1 _332_ (
  .A(_095_),
  .B1(_014_),
  .B2(_058_),
  .ZN(_091_)
);

NAND2_X1 _333_ (
  .A1(_090_),
  .A2(_091_),
  .ZN(_092_)
);

AOI21_X2 _334_ (
  .A(_085_),
  .B1(_089_),
  .B2(_092_),
  .ZN(_007_)
);

NAND2_X1 _335_ (
  .A1(_014_),
  .A2(_020_),
  .ZN(_093_)
);

MUX2_X1 _336_ (
  .A(\coef[30] ),
  .B(_093_),
  .S(_122_),
  .Z(_008_)
);

HA_X1 _337_ (
  .A(_163_),
  .B(_164_),
  .CO(_165_),
  .S(_166_)
);

HA_X1 _338_ (
  .A(_163_),
  .B(_164_),
  .CO(_167_),
  .S(_168_)
);

HA_X1 _339_ (
  .A(_163_),
  .B(x[1]),
  .CO(_169_),
  .S(_170_)
);

HA_X1 _340_ (
  .A(_163_),
  .B(x[1]),
  .CO(_171_),
  .S(_172_)
);

HA_X1 _341_ (
  .A(x[0]),
  .B(_164_),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _342_ (
  .A(x[0]),
  .B(_164_),
  .CO(_175_),
  .S(_176_)
);

HA_X1 _343_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_177_),
  .S(_178_)
);

HA_X1 _344_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_179_),
  .S(_180_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_162_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_161_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_160_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_159_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_158_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_157_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_156_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_155_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_154_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$5778094f610ca183dd46956f589e4ea513d2316c\dctu

module \$paramod$2da196d8114b669d4bb3858ca0a91434452576e0\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire \coef[10] ;
wire \coef[11] ;
wire \coef[13] ;
wire \coef[15] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

BUF_X4 _30_ (
  .A(y[2]),
  .Z(_04_)
);

INV_X4 _31_ (
  .A(_04_),
  .ZN(_05_)
);

NAND2_X2 _32_ (
  .A1(_05_),
  .A2(y[0]),
  .ZN(_06_)
);

INV_X1 _33_ (
  .A(y[0]),
  .ZN(_07_)
);

NAND2_X1 _34_ (
  .A1(_07_),
  .A2(_04_),
  .ZN(_08_)
);

BUF_X4 _35_ (
  .A(ena),
  .Z(_09_)
);

NAND3_X1 _36_ (
  .A1(_06_),
  .A2(_08_),
  .A3(_09_),
  .ZN(_10_)
);

INV_X2 _37_ (
  .A(_09_),
  .ZN(_11_)
);

NAND2_X1 _38_ (
  .A1(_11_),
  .A2(\coef[11] ),
  .ZN(_12_)
);

NAND2_X1 _39_ (
  .A1(_10_),
  .A2(_12_),
  .ZN(_00_)
);

NAND2_X2 _40_ (
  .A1(_05_),
  .A2(y[1]),
  .ZN(_13_)
);

INV_X1 _41_ (
  .A(y[1]),
  .ZN(_14_)
);

NAND2_X1 _42_ (
  .A1(_14_),
  .A2(_04_),
  .ZN(_15_)
);

NAND3_X1 _43_ (
  .A1(_13_),
  .A2(_15_),
  .A3(_09_),
  .ZN(_16_)
);

NAND2_X1 _44_ (
  .A1(_11_),
  .A2(\coef[13] ),
  .ZN(_17_)
);

NAND2_X1 _45_ (
  .A1(_16_),
  .A2(_17_),
  .ZN(_01_)
);

NAND2_X1 _46_ (
  .A1(_11_),
  .A2(\coef[10] ),
  .ZN(_18_)
);

NAND2_X1 _47_ (
  .A1(_04_),
  .A2(y[1]),
  .ZN(_19_)
);

NAND2_X1 _48_ (
  .A1(_19_),
  .A2(_09_),
  .ZN(_20_)
);

NOR2_X1 _49_ (
  .A1(_04_),
  .A2(y[1]),
  .ZN(_21_)
);

OAI21_X2 _50_ (
  .A(_18_),
  .B1(_20_),
  .B2(_21_),
  .ZN(_02_)
);

NAND2_X1 _51_ (
  .A1(_11_),
  .A2(\coef[15] ),
  .ZN(_22_)
);

NAND2_X1 _52_ (
  .A1(_04_),
  .A2(y[0]),
  .ZN(_23_)
);

NAND2_X1 _53_ (
  .A1(_23_),
  .A2(_09_),
  .ZN(_24_)
);

NOR2_X1 _54_ (
  .A1(_04_),
  .A2(y[0]),
  .ZN(_25_)
);

OAI21_X2 _55_ (
  .A(_22_),
  .B1(_24_),
  .B2(_25_),
  .ZN(_03_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[11] ),
  .QN(_29_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_01_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_28_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_02_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_27_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_03_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_26_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[15] , \coef[15] , \coef[10] , \coef[13] , \coef[10] , \coef[15] , \coef[15] , \coef[11] , \coef[10] , \coef[11] , \coef[15] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$2da196d8114b669d4bb3858ca0a91434452576e0\dctu

module \$paramod$696f85e1ea63d2b5ad7171a625fd3b51a665057d\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _185_ (
  .A(x[0]),
  .ZN(_167_)
);

INV_X1 _186_ (
  .A(x[1]),
  .ZN(_168_)
);

BUF_X8 _187_ (
  .A(x[2]),
  .Z(_098_)
);

INV_X8 _188_ (
  .A(_098_),
  .ZN(_099_)
);

BUF_X16 _189_ (
  .A(_099_),
  .Z(_100_)
);

INV_X1 _190_ (
  .A(_179_),
  .ZN(_101_)
);

NAND2_X4 _191_ (
  .A1(_100_),
  .A2(_101_),
  .ZN(_102_)
);

NAND2_X1 _192_ (
  .A1(_098_),
  .A2(_173_),
  .ZN(_103_)
);

NAND2_X2 _193_ (
  .A1(_102_),
  .A2(_103_),
  .ZN(_104_)
);

BUF_X4 _194_ (
  .A(y[0]),
  .Z(_105_)
);

BUF_X4 _195_ (
  .A(_105_),
  .Z(_106_)
);

NAND2_X2 _196_ (
  .A1(_104_),
  .A2(_106_),
  .ZN(_107_)
);

INV_X1 _197_ (
  .A(_170_),
  .ZN(_108_)
);

NAND2_X4 _198_ (
  .A1(_100_),
  .A2(_108_),
  .ZN(_109_)
);

NAND2_X1 _199_ (
  .A1(_098_),
  .A2(_170_),
  .ZN(_110_)
);

NAND2_X4 _200_ (
  .A1(_109_),
  .A2(_110_),
  .ZN(_111_)
);

INV_X4 _201_ (
  .A(_105_),
  .ZN(_112_)
);

BUF_X4 _202_ (
  .A(_112_),
  .Z(_113_)
);

NAND2_X4 _203_ (
  .A1(_111_),
  .A2(_113_),
  .ZN(_114_)
);

BUF_X2 _204_ (
  .A(y[1]),
  .Z(_115_)
);

CLKBUF_X3 _205_ (
  .A(_115_),
  .Z(_116_)
);

NAND3_X1 _206_ (
  .A1(_107_),
  .A2(_114_),
  .A3(_116_),
  .ZN(_117_)
);

BUF_X2 _207_ (
  .A(y[2]),
  .Z(_118_)
);

INV_X1 _208_ (
  .A(_169_),
  .ZN(_119_)
);

NAND2_X2 _209_ (
  .A1(_099_),
  .A2(_119_),
  .ZN(_120_)
);

NAND2_X1 _210_ (
  .A1(_098_),
  .A2(_183_),
  .ZN(_121_)
);

NAND3_X1 _211_ (
  .A1(_120_),
  .A2(_113_),
  .A3(_121_),
  .ZN(_122_)
);

INV_X1 _212_ (
  .A(_115_),
  .ZN(_123_)
);

BUF_X4 _213_ (
  .A(_123_),
  .Z(_124_)
);

NAND2_X1 _214_ (
  .A1(x[1]),
  .A2(_105_),
  .ZN(_125_)
);

NAND3_X1 _215_ (
  .A1(_122_),
  .A2(_124_),
  .A3(_125_),
  .ZN(_126_)
);

NAND3_X1 _216_ (
  .A1(_117_),
  .A2(_118_),
  .A3(_126_),
  .ZN(_127_)
);

NAND3_X2 _217_ (
  .A1(_109_),
  .A2(_106_),
  .A3(_110_),
  .ZN(_128_)
);

INV_X1 _218_ (
  .A(_177_),
  .ZN(_129_)
);

NAND2_X4 _219_ (
  .A1(_100_),
  .A2(_129_),
  .ZN(_130_)
);

NAND2_X1 _220_ (
  .A1(_098_),
  .A2(_175_),
  .ZN(_131_)
);

NAND3_X2 _221_ (
  .A1(_130_),
  .A2(_112_),
  .A3(_131_),
  .ZN(_132_)
);

NAND3_X1 _222_ (
  .A1(_128_),
  .A2(_132_),
  .A3(_124_),
  .ZN(_133_)
);

AOI21_X2 _223_ (
  .A(_123_),
  .B1(_113_),
  .B2(_168_),
  .ZN(_134_)
);

INV_X1 _224_ (
  .A(_171_),
  .ZN(_135_)
);

NAND2_X4 _225_ (
  .A1(_100_),
  .A2(_135_),
  .ZN(_136_)
);

NAND2_X1 _226_ (
  .A1(_098_),
  .A2(_181_),
  .ZN(_137_)
);

NAND2_X2 _227_ (
  .A1(_136_),
  .A2(_137_),
  .ZN(_138_)
);

INV_X1 _228_ (
  .A(_138_),
  .ZN(_139_)
);

OAI21_X1 _229_ (
  .A(_134_),
  .B1(_139_),
  .B2(_113_),
  .ZN(_140_)
);

INV_X2 _230_ (
  .A(_118_),
  .ZN(_141_)
);

NAND3_X1 _231_ (
  .A1(_133_),
  .A2(_140_),
  .A3(_141_),
  .ZN(_142_)
);

BUF_X4 _232_ (
  .A(ena),
  .Z(_143_)
);

NAND3_X1 _233_ (
  .A1(_127_),
  .A2(_142_),
  .A3(_143_),
  .ZN(_144_)
);

INV_X2 _234_ (
  .A(_143_),
  .ZN(_145_)
);

NAND2_X1 _235_ (
  .A1(_145_),
  .A2(\coef[21] ),
  .ZN(_146_)
);

NAND2_X1 _236_ (
  .A1(_144_),
  .A2(_146_),
  .ZN(_000_)
);

NAND2_X2 _237_ (
  .A1(_120_),
  .A2(_121_),
  .ZN(_147_)
);

NAND3_X1 _238_ (
  .A1(_147_),
  .A2(_106_),
  .A3(_124_),
  .ZN(_148_)
);

NAND2_X4 _239_ (
  .A1(_130_),
  .A2(_131_),
  .ZN(_149_)
);

NAND3_X1 _240_ (
  .A1(_149_),
  .A2(_106_),
  .A3(_116_),
  .ZN(_150_)
);

NAND4_X1 _241_ (
  .A1(_148_),
  .A2(_150_),
  .A3(_118_),
  .A4(_114_),
  .ZN(_151_)
);

NAND2_X1 _242_ (
  .A1(_138_),
  .A2(_115_),
  .ZN(_152_)
);

NAND2_X1 _243_ (
  .A1(_104_),
  .A2(_124_),
  .ZN(_153_)
);

NAND3_X1 _244_ (
  .A1(_152_),
  .A2(_153_),
  .A3(_113_),
  .ZN(_154_)
);

NAND3_X1 _245_ (
  .A1(_154_),
  .A2(_141_),
  .A3(_128_),
  .ZN(_155_)
);

NAND3_X1 _246_ (
  .A1(_151_),
  .A2(_155_),
  .A3(_143_),
  .ZN(_156_)
);

NAND2_X1 _247_ (
  .A1(_145_),
  .A2(\coef[23] ),
  .ZN(_157_)
);

NAND2_X1 _248_ (
  .A1(_156_),
  .A2(_157_),
  .ZN(_001_)
);

NOR2_X1 _249_ (
  .A1(_143_),
  .A2(\coef[24] ),
  .ZN(_009_)
);

AOI21_X1 _250_ (
  .A(_115_),
  .B1(_113_),
  .B2(x[0]),
  .ZN(_010_)
);

AOI21_X1 _251_ (
  .A(_118_),
  .B1(_128_),
  .B2(_010_),
  .ZN(_011_)
);

NAND2_X1 _252_ (
  .A1(_147_),
  .A2(_105_),
  .ZN(_012_)
);

NAND2_X4 _253_ (
  .A1(_100_),
  .A2(_181_),
  .ZN(_013_)
);

NAND2_X1 _254_ (
  .A1(_135_),
  .A2(_098_),
  .ZN(_014_)
);

NAND3_X2 _255_ (
  .A1(_013_),
  .A2(_014_),
  .A3(_112_),
  .ZN(_015_)
);

NAND3_X1 _256_ (
  .A1(_012_),
  .A2(_015_),
  .A3(_115_),
  .ZN(_016_)
);

AOI21_X1 _257_ (
  .A(_145_),
  .B1(_011_),
  .B2(_016_),
  .ZN(_017_)
);

NAND3_X2 _258_ (
  .A1(_136_),
  .A2(_112_),
  .A3(_137_),
  .ZN(_018_)
);

INV_X1 _259_ (
  .A(_183_),
  .ZN(_019_)
);

NAND2_X4 _260_ (
  .A1(_100_),
  .A2(_019_),
  .ZN(_020_)
);

NAND2_X1 _261_ (
  .A1(_098_),
  .A2(_169_),
  .ZN(_021_)
);

NAND3_X1 _262_ (
  .A1(_020_),
  .A2(_105_),
  .A3(_021_),
  .ZN(_022_)
);

NAND3_X1 _263_ (
  .A1(_018_),
  .A2(_022_),
  .A3(_124_),
  .ZN(_023_)
);

NOR2_X1 _264_ (
  .A1(_112_),
  .A2(x[0]),
  .ZN(_024_)
);

INV_X1 _265_ (
  .A(_024_),
  .ZN(_025_)
);

NAND3_X1 _266_ (
  .A1(_114_),
  .A2(_116_),
  .A3(_025_),
  .ZN(_026_)
);

NAND3_X1 _267_ (
  .A1(_023_),
  .A2(_026_),
  .A3(_118_),
  .ZN(_027_)
);

AOI21_X2 _268_ (
  .A(_009_),
  .B1(_017_),
  .B2(_027_),
  .ZN(_002_)
);

NOR2_X1 _269_ (
  .A1(_143_),
  .A2(\coef[10] ),
  .ZN(_028_)
);

NAND2_X1 _270_ (
  .A1(_100_),
  .A2(_106_),
  .ZN(_029_)
);

AOI21_X1 _271_ (
  .A(_141_),
  .B1(_010_),
  .B2(_029_),
  .ZN(_030_)
);

NAND2_X1 _272_ (
  .A1(_111_),
  .A2(_106_),
  .ZN(_031_)
);

NAND2_X1 _273_ (
  .A1(_031_),
  .A2(_134_),
  .ZN(_032_)
);

AOI21_X1 _274_ (
  .A(_145_),
  .B1(_030_),
  .B2(_032_),
  .ZN(_033_)
);

NAND3_X2 _275_ (
  .A1(_109_),
  .A2(_113_),
  .A3(_110_),
  .ZN(_034_)
);

NAND2_X1 _276_ (
  .A1(_125_),
  .A2(_123_),
  .ZN(_035_)
);

INV_X1 _277_ (
  .A(_035_),
  .ZN(_036_)
);

AOI21_X2 _278_ (
  .A(_118_),
  .B1(_034_),
  .B2(_036_),
  .ZN(_037_)
);

NOR2_X1 _279_ (
  .A1(_100_),
  .A2(_105_),
  .ZN(_038_)
);

INV_X1 _280_ (
  .A(_038_),
  .ZN(_039_)
);

NAND3_X1 _281_ (
  .A1(_025_),
  .A2(_039_),
  .A3(_116_),
  .ZN(_040_)
);

NAND2_X1 _282_ (
  .A1(_037_),
  .A2(_040_),
  .ZN(_041_)
);

AOI21_X2 _283_ (
  .A(_028_),
  .B1(_033_),
  .B2(_041_),
  .ZN(_003_)
);

NAND3_X1 _284_ (
  .A1(_107_),
  .A2(_132_),
  .A3(_124_),
  .ZN(_042_)
);

NAND3_X1 _285_ (
  .A1(_042_),
  .A2(_032_),
  .A3(_118_),
  .ZN(_043_)
);

NAND3_X1 _286_ (
  .A1(_107_),
  .A2(_132_),
  .A3(_116_),
  .ZN(_044_)
);

NAND2_X1 _287_ (
  .A1(_037_),
  .A2(_044_),
  .ZN(_045_)
);

NAND3_X1 _288_ (
  .A1(_043_),
  .A2(_143_),
  .A3(_045_),
  .ZN(_046_)
);

NAND2_X1 _289_ (
  .A1(_145_),
  .A2(\coef[26] ),
  .ZN(_047_)
);

NAND2_X1 _290_ (
  .A1(_046_),
  .A2(_047_),
  .ZN(_004_)
);

NOR2_X1 _291_ (
  .A1(_143_),
  .A2(\coef[13] ),
  .ZN(_048_)
);

NAND2_X4 _292_ (
  .A1(_100_),
  .A2(_173_),
  .ZN(_049_)
);

NAND2_X1 _293_ (
  .A1(_101_),
  .A2(_098_),
  .ZN(_050_)
);

NAND2_X2 _294_ (
  .A1(_049_),
  .A2(_050_),
  .ZN(_051_)
);

NAND2_X2 _295_ (
  .A1(_051_),
  .A2(_106_),
  .ZN(_052_)
);

NAND3_X1 _296_ (
  .A1(_052_),
  .A2(_116_),
  .A3(_039_),
  .ZN(_053_)
);

INV_X1 _297_ (
  .A(_053_),
  .ZN(_054_)
);

NAND3_X1 _298_ (
  .A1(_020_),
  .A2(_113_),
  .A3(_021_),
  .ZN(_055_)
);

AOI21_X1 _299_ (
  .A(_116_),
  .B1(_055_),
  .B2(_025_),
  .ZN(_056_)
);

OAI21_X1 _300_ (
  .A(_141_),
  .B1(_054_),
  .B2(_056_),
  .ZN(_057_)
);

NAND3_X1 _301_ (
  .A1(_013_),
  .A2(_014_),
  .A3(_106_),
  .ZN(_058_)
);

NAND2_X1 _302_ (
  .A1(_112_),
  .A2(x[0]),
  .ZN(_059_)
);

NAND2_X1 _303_ (
  .A1(_059_),
  .A2(_115_),
  .ZN(_060_)
);

INV_X1 _304_ (
  .A(_060_),
  .ZN(_061_)
);

AOI21_X1 _305_ (
  .A(_141_),
  .B1(_058_),
  .B2(_061_),
  .ZN(_062_)
);

INV_X1 _306_ (
  .A(_175_),
  .ZN(_063_)
);

NAND2_X4 _307_ (
  .A1(_100_),
  .A2(_063_),
  .ZN(_064_)
);

NAND2_X1 _308_ (
  .A1(_098_),
  .A2(_177_),
  .ZN(_065_)
);

NAND2_X2 _309_ (
  .A1(_064_),
  .A2(_065_),
  .ZN(_066_)
);

NAND2_X2 _310_ (
  .A1(_066_),
  .A2(_113_),
  .ZN(_067_)
);

NAND2_X2 _311_ (
  .A1(_067_),
  .A2(_029_),
  .ZN(_068_)
);

NAND2_X1 _312_ (
  .A1(_068_),
  .A2(_124_),
  .ZN(_069_)
);

AOI21_X1 _313_ (
  .A(_145_),
  .B1(_062_),
  .B2(_069_),
  .ZN(_070_)
);

AOI21_X1 _314_ (
  .A(_048_),
  .B1(_057_),
  .B2(_070_),
  .ZN(_005_)
);

NAND2_X1 _315_ (
  .A1(_149_),
  .A2(_113_),
  .ZN(_071_)
);

NAND3_X1 _316_ (
  .A1(_064_),
  .A2(_106_),
  .A3(_065_),
  .ZN(_072_)
);

NAND3_X1 _317_ (
  .A1(_071_),
  .A2(_072_),
  .A3(_116_),
  .ZN(_073_)
);

NAND3_X1 _318_ (
  .A1(_023_),
  .A2(_073_),
  .A3(_118_),
  .ZN(_074_)
);

NAND3_X1 _319_ (
  .A1(_049_),
  .A2(_050_),
  .A3(_112_),
  .ZN(_075_)
);

NAND3_X1 _320_ (
  .A1(_102_),
  .A2(_105_),
  .A3(_103_),
  .ZN(_076_)
);

NAND3_X1 _321_ (
  .A1(_075_),
  .A2(_076_),
  .A3(_124_),
  .ZN(_077_)
);

NAND3_X1 _322_ (
  .A1(_016_),
  .A2(_077_),
  .A3(_141_),
  .ZN(_078_)
);

NAND2_X1 _323_ (
  .A1(_074_),
  .A2(_078_),
  .ZN(_079_)
);

NAND2_X1 _324_ (
  .A1(_079_),
  .A2(_143_),
  .ZN(_080_)
);

NAND2_X1 _325_ (
  .A1(_145_),
  .A2(\coef[28] ),
  .ZN(_081_)
);

NAND2_X1 _326_ (
  .A1(_080_),
  .A2(_081_),
  .ZN(_006_)
);

NAND2_X1 _327_ (
  .A1(_012_),
  .A2(_059_),
  .ZN(_082_)
);

NAND2_X1 _328_ (
  .A1(_082_),
  .A2(_116_),
  .ZN(_083_)
);

NOR2_X1 _329_ (
  .A1(_168_),
  .A2(_105_),
  .ZN(_084_)
);

INV_X1 _330_ (
  .A(_084_),
  .ZN(_085_)
);

NAND3_X1 _331_ (
  .A1(_052_),
  .A2(_124_),
  .A3(_085_),
  .ZN(_086_)
);

NAND3_X1 _332_ (
  .A1(_083_),
  .A2(_086_),
  .A3(_141_),
  .ZN(_087_)
);

NAND2_X1 _333_ (
  .A1(_018_),
  .A2(_025_),
  .ZN(_088_)
);

NAND2_X1 _334_ (
  .A1(_088_),
  .A2(_124_),
  .ZN(_089_)
);

NAND2_X1 _335_ (
  .A1(_168_),
  .A2(_106_),
  .ZN(_090_)
);

NAND3_X1 _336_ (
  .A1(_067_),
  .A2(_116_),
  .A3(_090_),
  .ZN(_091_)
);

NAND3_X1 _337_ (
  .A1(_089_),
  .A2(_091_),
  .A3(_118_),
  .ZN(_092_)
);

NAND3_X1 _338_ (
  .A1(_087_),
  .A2(_092_),
  .A3(_143_),
  .ZN(_093_)
);

NAND2_X1 _339_ (
  .A1(_145_),
  .A2(\coef[29] ),
  .ZN(_094_)
);

NAND2_X1 _340_ (
  .A1(_093_),
  .A2(_094_),
  .ZN(_007_)
);

NOR2_X1 _341_ (
  .A1(_143_),
  .A2(\coef[30] ),
  .ZN(_095_)
);

AOI21_X1 _342_ (
  .A(_145_),
  .B1(_147_),
  .B2(_141_),
  .ZN(_096_)
);

NAND2_X1 _343_ (
  .A1(_139_),
  .A2(_118_),
  .ZN(_097_)
);

AOI21_X1 _344_ (
  .A(_095_),
  .B1(_096_),
  .B2(_097_),
  .ZN(_008_)
);

HA_X1 _345_ (
  .A(_167_),
  .B(_168_),
  .CO(_169_),
  .S(_170_)
);

HA_X1 _346_ (
  .A(_167_),
  .B(_168_),
  .CO(_171_),
  .S(_172_)
);

HA_X1 _347_ (
  .A(_167_),
  .B(x[1]),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _348_ (
  .A(_167_),
  .B(x[1]),
  .CO(_175_),
  .S(_176_)
);

HA_X1 _349_ (
  .A(x[0]),
  .B(_168_),
  .CO(_177_),
  .S(_178_)
);

HA_X1 _350_ (
  .A(x[0]),
  .B(_168_),
  .CO(_179_),
  .S(_180_)
);

HA_X1 _351_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_181_),
  .S(_182_)
);

HA_X1 _352_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_183_),
  .S(_184_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_166_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_165_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_164_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_163_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_162_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_161_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_160_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_159_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_158_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$696f85e1ea63d2b5ad7171a625fd3b51a665057d\dctu

module \$paramod$6be19b0824fdb8c44e931702b04949b1ae101a34\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire \coef[10] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _068_ (
  .A(x[0]),
  .ZN(_058_)
);

INV_X1 _069_ (
  .A(x[1]),
  .ZN(_059_)
);

BUF_X8 _070_ (
  .A(y[0]),
  .Z(_003_)
);

NAND2_X1 _071_ (
  .A1(_003_),
  .A2(_066_),
  .ZN(_004_)
);

INV_X1 _072_ (
  .A(_062_),
  .ZN(_005_)
);

OAI21_X1 _073_ (
  .A(_004_),
  .B1(_003_),
  .B2(_005_),
  .ZN(_006_)
);

NOR2_X1 _074_ (
  .A1(_006_),
  .A2(y[1]),
  .ZN(_007_)
);

NOR2_X2 _075_ (
  .A1(_007_),
  .A2(y[2]),
  .ZN(_008_)
);

INV_X8 _076_ (
  .A(_003_),
  .ZN(_009_)
);

BUF_X4 _077_ (
  .A(x[2]),
  .Z(_010_)
);

NAND2_X2 _078_ (
  .A1(_009_),
  .A2(_010_),
  .ZN(_011_)
);

NAND2_X4 _079_ (
  .A1(_009_),
  .A2(_061_),
  .ZN(_012_)
);

NAND2_X4 _080_ (
  .A1(_011_),
  .A2(_012_),
  .ZN(_013_)
);

INV_X2 _081_ (
  .A(_010_),
  .ZN(_014_)
);

OAI21_X2 _082_ (
  .A(_013_),
  .B1(_066_),
  .B2(_014_),
  .ZN(_015_)
);

NAND3_X1 _083_ (
  .A1(_003_),
  .A2(_062_),
  .A3(_010_),
  .ZN(_016_)
);

NAND2_X1 _084_ (
  .A1(_016_),
  .A2(y[1]),
  .ZN(_017_)
);

INV_X1 _085_ (
  .A(_017_),
  .ZN(_018_)
);

NAND2_X2 _086_ (
  .A1(_015_),
  .A2(_018_),
  .ZN(_019_)
);

NAND2_X2 _087_ (
  .A1(_008_),
  .A2(_019_),
  .ZN(_020_)
);

NAND2_X1 _088_ (
  .A1(_005_),
  .A2(_010_),
  .ZN(_021_)
);

NAND2_X1 _089_ (
  .A1(_014_),
  .A2(_061_),
  .ZN(_022_)
);

NAND3_X1 _090_ (
  .A1(_021_),
  .A2(_022_),
  .A3(_009_),
  .ZN(_023_)
);

INV_X2 _091_ (
  .A(y[1]),
  .ZN(_024_)
);

NAND3_X1 _092_ (
  .A1(_003_),
  .A2(_066_),
  .A3(_010_),
  .ZN(_025_)
);

NAND3_X1 _093_ (
  .A1(_023_),
  .A2(_024_),
  .A3(_025_),
  .ZN(_026_)
);

NAND2_X2 _094_ (
  .A1(_012_),
  .A2(y[1]),
  .ZN(_027_)
);

AND2_X2 _095_ (
  .A1(_027_),
  .A2(y[2]),
  .ZN(_028_)
);

NAND2_X1 _096_ (
  .A1(_026_),
  .A2(_028_),
  .ZN(_029_)
);

NAND2_X2 _097_ (
  .A1(_020_),
  .A2(_029_),
  .ZN(_030_)
);

BUF_X1 _098_ (
  .A(ena),
  .Z(_031_)
);

NAND2_X2 _099_ (
  .A1(_030_),
  .A2(_031_),
  .ZN(_032_)
);

INV_X1 _100_ (
  .A(_031_),
  .ZN(_033_)
);

NAND2_X1 _101_ (
  .A1(_033_),
  .A2(\coef[10] ),
  .ZN(_034_)
);

NAND2_X2 _102_ (
  .A1(_032_),
  .A2(_034_),
  .ZN(_000_)
);

NOR2_X1 _103_ (
  .A1(_031_),
  .A2(\coef[29] ),
  .ZN(_035_)
);

NAND2_X1 _104_ (
  .A1(_010_),
  .A2(_060_),
  .ZN(_036_)
);

NAND2_X2 _105_ (
  .A1(_013_),
  .A2(_036_),
  .ZN(_037_)
);

NAND2_X1 _106_ (
  .A1(_010_),
  .A2(_064_),
  .ZN(_038_)
);

NAND2_X1 _107_ (
  .A1(_038_),
  .A2(_003_),
  .ZN(_039_)
);

NAND2_X2 _108_ (
  .A1(_037_),
  .A2(_039_),
  .ZN(_040_)
);

NAND2_X2 _109_ (
  .A1(_040_),
  .A2(_024_),
  .ZN(_041_)
);

NAND2_X2 _110_ (
  .A1(_041_),
  .A2(_027_),
  .ZN(_042_)
);

NAND2_X2 _111_ (
  .A1(_042_),
  .A2(y[2]),
  .ZN(_043_)
);

NAND2_X1 _112_ (
  .A1(_009_),
  .A2(_060_),
  .ZN(_044_)
);

NAND2_X1 _113_ (
  .A1(_003_),
  .A2(_064_),
  .ZN(_045_)
);

NAND2_X1 _114_ (
  .A1(_044_),
  .A2(_045_),
  .ZN(_046_)
);

AOI21_X1 _115_ (
  .A(y[2]),
  .B1(_046_),
  .B2(_024_),
  .ZN(_047_)
);

AOI21_X1 _116_ (
  .A(_024_),
  .B1(_036_),
  .B2(_003_),
  .ZN(_048_)
);

NAND3_X1 _117_ (
  .A1(_022_),
  .A2(_038_),
  .A3(_009_),
  .ZN(_049_)
);

NAND2_X1 _118_ (
  .A1(_048_),
  .A2(_049_),
  .ZN(_050_)
);

AOI21_X1 _119_ (
  .A(_033_),
  .B1(_047_),
  .B2(_050_),
  .ZN(_051_)
);

AOI21_X2 _120_ (
  .A(_035_),
  .B1(_043_),
  .B2(_051_),
  .ZN(_001_)
);

NOR2_X1 _121_ (
  .A1(_031_),
  .A2(\coef[30] ),
  .ZN(_052_)
);

XNOR2_X1 _122_ (
  .A(_003_),
  .B(_061_),
  .ZN(_053_)
);

XNOR2_X1 _123_ (
  .A(_053_),
  .B(_024_),
  .ZN(_054_)
);

AOI21_X1 _124_ (
  .A(_052_),
  .B1(_054_),
  .B2(_031_),
  .ZN(_002_)
);

HA_X1 _125_ (
  .A(_058_),
  .B(_059_),
  .CO(_060_),
  .S(_061_)
);

HA_X1 _126_ (
  .A(_058_),
  .B(_059_),
  .CO(_062_),
  .S(_063_)
);

HA_X1 _127_ (
  .A(_058_),
  .B(x[1]),
  .CO(_064_),
  .S(_065_)
);

HA_X1 _128_ (
  .A(_058_),
  .B(x[1]),
  .CO(_066_),
  .S(_067_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_057_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_056_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_055_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[10] , \coef[10] , \coef[10] , \coef[10] , \coef[10] , \coef[10] , \coef[10] , \coef[10] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$6be19b0824fdb8c44e931702b04949b1ae101a34\dctu

module \$paramod$785fe1ea8cdf428cbeb2f89081ee68c33feb7da2\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _202_ (
  .A(x[1]),
  .ZN(_185_)
);

INV_X1 _203_ (
  .A(x[0]),
  .ZN(_184_)
);

INV_X2 _204_ (
  .A(x[2]),
  .ZN(_115_)
);

INV_X1 _205_ (
  .A(_198_),
  .ZN(_116_)
);

NAND2_X1 _206_ (
  .A1(_115_),
  .A2(_116_),
  .ZN(_117_)
);

NAND2_X1 _207_ (
  .A1(x[2]),
  .A2(_188_),
  .ZN(_118_)
);

NAND2_X1 _208_ (
  .A1(_117_),
  .A2(_118_),
  .ZN(_119_)
);

BUF_X4 _209_ (
  .A(y[0]),
  .Z(_120_)
);

BUF_X4 _210_ (
  .A(_120_),
  .Z(_121_)
);

NAND2_X1 _211_ (
  .A1(_119_),
  .A2(_121_),
  .ZN(_122_)
);

BUF_X2 _212_ (
  .A(y[1]),
  .Z(_123_)
);

INV_X2 _213_ (
  .A(_123_),
  .ZN(_124_)
);

INV_X2 _214_ (
  .A(_120_),
  .ZN(_125_)
);

BUF_X8 _215_ (
  .A(_125_),
  .Z(_126_)
);

AOI21_X2 _216_ (
  .A(_124_),
  .B1(_184_),
  .B2(_126_),
  .ZN(_127_)
);

NAND2_X1 _217_ (
  .A1(_122_),
  .A2(_127_),
  .ZN(_128_)
);

BUF_X8 _218_ (
  .A(_115_),
  .Z(_129_)
);

NAND2_X2 _219_ (
  .A1(_129_),
  .A2(_190_),
  .ZN(_130_)
);

INV_X1 _220_ (
  .A(_196_),
  .ZN(_131_)
);

BUF_X4 _221_ (
  .A(x[2]),
  .Z(_132_)
);

NAND2_X1 _222_ (
  .A1(_131_),
  .A2(_132_),
  .ZN(_133_)
);

NAND3_X1 _223_ (
  .A1(_130_),
  .A2(_133_),
  .A3(_126_),
  .ZN(_134_)
);

NAND2_X1 _224_ (
  .A1(_132_),
  .A2(_120_),
  .ZN(_135_)
);

NAND2_X1 _225_ (
  .A1(_135_),
  .A2(_124_),
  .ZN(_136_)
);

INV_X1 _226_ (
  .A(_136_),
  .ZN(_137_)
);

NAND2_X1 _227_ (
  .A1(_134_),
  .A2(_137_),
  .ZN(_138_)
);

BUF_X2 _228_ (
  .A(y[2]),
  .Z(_139_)
);

INV_X1 _229_ (
  .A(_139_),
  .ZN(_140_)
);

NAND3_X1 _230_ (
  .A1(_128_),
  .A2(_138_),
  .A3(_140_),
  .ZN(_141_)
);

INV_X1 _231_ (
  .A(_192_),
  .ZN(_142_)
);

NAND2_X1 _232_ (
  .A1(_129_),
  .A2(_142_),
  .ZN(_143_)
);

NAND2_X1 _233_ (
  .A1(_132_),
  .A2(_194_),
  .ZN(_144_)
);

NAND3_X1 _234_ (
  .A1(_143_),
  .A2(_121_),
  .A3(_144_),
  .ZN(_145_)
);

AOI21_X1 _235_ (
  .A(_124_),
  .B1(_126_),
  .B2(_129_),
  .ZN(_146_)
);

NAND2_X1 _236_ (
  .A1(_145_),
  .A2(_146_),
  .ZN(_147_)
);

INV_X1 _237_ (
  .A(_200_),
  .ZN(_148_)
);

NAND2_X1 _238_ (
  .A1(_129_),
  .A2(_148_),
  .ZN(_149_)
);

NAND2_X1 _239_ (
  .A1(_132_),
  .A2(_186_),
  .ZN(_150_)
);

NAND3_X1 _240_ (
  .A1(_149_),
  .A2(_126_),
  .A3(_150_),
  .ZN(_151_)
);

NAND2_X1 _241_ (
  .A1(_120_),
  .A2(x[0]),
  .ZN(_152_)
);

NAND2_X1 _242_ (
  .A1(_152_),
  .A2(_124_),
  .ZN(_153_)
);

INV_X1 _243_ (
  .A(_153_),
  .ZN(_154_)
);

NAND2_X1 _244_ (
  .A1(_151_),
  .A2(_154_),
  .ZN(_155_)
);

NAND3_X1 _245_ (
  .A1(_147_),
  .A2(_155_),
  .A3(_139_),
  .ZN(_156_)
);

BUF_X1 _246_ (
  .A(ena),
  .Z(_157_)
);

NAND3_X1 _247_ (
  .A1(_141_),
  .A2(_156_),
  .A3(_157_),
  .ZN(_158_)
);

OR2_X1 _248_ (
  .A1(_157_),
  .A2(\coef[21] ),
  .ZN(_159_)
);

AND2_X2 _249_ (
  .A1(_158_),
  .A2(_159_),
  .ZN(_000_)
);

NOR2_X1 _250_ (
  .A1(_157_),
  .A2(\coef[23] ),
  .ZN(_160_)
);

OAI21_X1 _251_ (
  .A(_152_),
  .B1(_129_),
  .B2(_121_),
  .ZN(_161_)
);

BUF_X2 _252_ (
  .A(_124_),
  .Z(_162_)
);

OAI21_X1 _253_ (
  .A(_139_),
  .B1(_161_),
  .B2(_162_),
  .ZN(_163_)
);

INV_X1 _254_ (
  .A(_163_),
  .ZN(_164_)
);

BUF_X2 _255_ (
  .A(_123_),
  .Z(_165_)
);

OAI21_X1 _256_ (
  .A(_164_),
  .B1(_165_),
  .B2(_119_),
  .ZN(_166_)
);

INV_X1 _257_ (
  .A(ena),
  .ZN(_167_)
);

OAI21_X1 _258_ (
  .A(_135_),
  .B1(_121_),
  .B2(_184_),
  .ZN(_168_)
);

AOI21_X1 _259_ (
  .A(_139_),
  .B1(_168_),
  .B2(_162_),
  .ZN(_169_)
);

NAND2_X1 _260_ (
  .A1(_129_),
  .A2(_200_),
  .ZN(_170_)
);

INV_X1 _261_ (
  .A(_186_),
  .ZN(_171_)
);

NAND2_X1 _262_ (
  .A1(_171_),
  .A2(_132_),
  .ZN(_172_)
);

NAND3_X1 _263_ (
  .A1(_170_),
  .A2(_172_),
  .A3(_165_),
  .ZN(_173_)
);

AOI21_X1 _264_ (
  .A(_167_),
  .B1(_169_),
  .B2(_173_),
  .ZN(_174_)
);

AOI21_X1 _265_ (
  .A(_160_),
  .B1(_166_),
  .B2(_174_),
  .ZN(_001_)
);

NAND3_X1 _266_ (
  .A1(_170_),
  .A2(_172_),
  .A3(_121_),
  .ZN(_009_)
);

AOI21_X1 _267_ (
  .A(_139_),
  .B1(_009_),
  .B2(_127_),
  .ZN(_010_)
);

INV_X1 _268_ (
  .A(_194_),
  .ZN(_011_)
);

NAND2_X1 _269_ (
  .A1(_115_),
  .A2(_011_),
  .ZN(_012_)
);

NAND2_X1 _270_ (
  .A1(_132_),
  .A2(_192_),
  .ZN(_013_)
);

NAND2_X1 _271_ (
  .A1(_012_),
  .A2(_013_),
  .ZN(_014_)
);

NAND2_X1 _272_ (
  .A1(_014_),
  .A2(_121_),
  .ZN(_015_)
);

NAND2_X1 _273_ (
  .A1(_125_),
  .A2(x[1]),
  .ZN(_016_)
);

NAND2_X1 _274_ (
  .A1(_015_),
  .A2(_016_),
  .ZN(_017_)
);

NAND2_X1 _275_ (
  .A1(_017_),
  .A2(_162_),
  .ZN(_018_)
);

NAND2_X1 _276_ (
  .A1(_010_),
  .A2(_018_),
  .ZN(_019_)
);

NAND3_X1 _277_ (
  .A1(_117_),
  .A2(_126_),
  .A3(_118_),
  .ZN(_020_)
);

AOI21_X1 _278_ (
  .A(_140_),
  .B1(_020_),
  .B2(_154_),
  .ZN(_021_)
);

NAND2_X4 _279_ (
  .A1(_129_),
  .A2(_131_),
  .ZN(_022_)
);

NAND2_X1 _280_ (
  .A1(_132_),
  .A2(_190_),
  .ZN(_023_)
);

NAND3_X2 _281_ (
  .A1(_022_),
  .A2(_126_),
  .A3(_023_),
  .ZN(_024_)
);

NAND2_X1 _282_ (
  .A1(_185_),
  .A2(_121_),
  .ZN(_025_)
);

NAND2_X1 _283_ (
  .A1(_024_),
  .A2(_025_),
  .ZN(_026_)
);

NAND2_X1 _284_ (
  .A1(_026_),
  .A2(_165_),
  .ZN(_027_)
);

NAND2_X1 _285_ (
  .A1(_021_),
  .A2(_027_),
  .ZN(_028_)
);

NAND3_X1 _286_ (
  .A1(_019_),
  .A2(_028_),
  .A3(_157_),
  .ZN(_029_)
);

NAND2_X1 _287_ (
  .A1(_167_),
  .A2(\coef[24] ),
  .ZN(_030_)
);

NAND2_X1 _288_ (
  .A1(_029_),
  .A2(_030_),
  .ZN(_002_)
);

NAND3_X1 _289_ (
  .A1(_143_),
  .A2(_126_),
  .A3(_144_),
  .ZN(_031_)
);

NOR2_X1 _290_ (
  .A1(_031_),
  .A2(_165_),
  .ZN(_032_)
);

NOR2_X1 _291_ (
  .A1(_125_),
  .A2(_123_),
  .ZN(_033_)
);

NAND3_X1 _292_ (
  .A1(_033_),
  .A2(_022_),
  .A3(_023_),
  .ZN(_034_)
);

NAND2_X1 _293_ (
  .A1(_034_),
  .A2(_139_),
  .ZN(_035_)
);

NOR2_X1 _294_ (
  .A1(_032_),
  .A2(_035_),
  .ZN(_036_)
);

NAND2_X1 _295_ (
  .A1(_129_),
  .A2(_171_),
  .ZN(_037_)
);

NAND2_X1 _296_ (
  .A1(_132_),
  .A2(_200_),
  .ZN(_038_)
);

NAND2_X1 _297_ (
  .A1(_037_),
  .A2(_038_),
  .ZN(_039_)
);

NAND2_X1 _298_ (
  .A1(_039_),
  .A2(_121_),
  .ZN(_040_)
);

NAND2_X1 _299_ (
  .A1(_040_),
  .A2(_151_),
  .ZN(_041_)
);

NAND2_X1 _300_ (
  .A1(_041_),
  .A2(_165_),
  .ZN(_042_)
);

NAND2_X1 _301_ (
  .A1(_036_),
  .A2(_042_),
  .ZN(_043_)
);

NAND3_X1 _302_ (
  .A1(_130_),
  .A2(_133_),
  .A3(_121_),
  .ZN(_044_)
);

NOR2_X1 _303_ (
  .A1(_044_),
  .A2(_124_),
  .ZN(_045_)
);

NOR2_X1 _304_ (
  .A1(_124_),
  .A2(_120_),
  .ZN(_046_)
);

NAND2_X1 _305_ (
  .A1(_014_),
  .A2(_046_),
  .ZN(_047_)
);

NAND2_X1 _306_ (
  .A1(_047_),
  .A2(_140_),
  .ZN(_048_)
);

NOR2_X1 _307_ (
  .A1(_045_),
  .A2(_048_),
  .ZN(_049_)
);

NAND2_X1 _308_ (
  .A1(_115_),
  .A2(_188_),
  .ZN(_050_)
);

NAND2_X1 _309_ (
  .A1(_116_),
  .A2(_132_),
  .ZN(_051_)
);

NAND2_X1 _310_ (
  .A1(_050_),
  .A2(_051_),
  .ZN(_052_)
);

NAND2_X1 _311_ (
  .A1(_052_),
  .A2(_126_),
  .ZN(_053_)
);

NAND2_X1 _312_ (
  .A1(_122_),
  .A2(_053_),
  .ZN(_054_)
);

NAND2_X1 _313_ (
  .A1(_054_),
  .A2(_162_),
  .ZN(_055_)
);

NAND2_X1 _314_ (
  .A1(_049_),
  .A2(_055_),
  .ZN(_056_)
);

NAND3_X1 _315_ (
  .A1(_043_),
  .A2(_056_),
  .A3(_157_),
  .ZN(_057_)
);

NAND2_X1 _316_ (
  .A1(_167_),
  .A2(\coef[10] ),
  .ZN(_058_)
);

NAND2_X1 _317_ (
  .A1(_057_),
  .A2(_058_),
  .ZN(_003_)
);

INV_X1 _318_ (
  .A(_145_),
  .ZN(_059_)
);

NOR2_X1 _319_ (
  .A1(_129_),
  .A2(_120_),
  .ZN(_060_)
);

OAI21_X1 _320_ (
  .A(_165_),
  .B1(_059_),
  .B2(_060_),
  .ZN(_061_)
);

NOR2_X1 _321_ (
  .A1(_060_),
  .A2(_165_),
  .ZN(_062_)
);

AOI21_X1 _322_ (
  .A(_139_),
  .B1(_009_),
  .B2(_062_),
  .ZN(_063_)
);

NAND2_X1 _323_ (
  .A1(_061_),
  .A2(_063_),
  .ZN(_064_)
);

NAND2_X1 _324_ (
  .A1(_129_),
  .A2(_120_),
  .ZN(_065_)
);

NAND2_X1 _325_ (
  .A1(_065_),
  .A2(_123_),
  .ZN(_066_)
);

INV_X1 _326_ (
  .A(_066_),
  .ZN(_067_)
);

AOI21_X1 _327_ (
  .A(_140_),
  .B1(_020_),
  .B2(_067_),
  .ZN(_068_)
);

NAND2_X1 _328_ (
  .A1(_134_),
  .A2(_065_),
  .ZN(_069_)
);

NAND2_X1 _329_ (
  .A1(_069_),
  .A2(_162_),
  .ZN(_070_)
);

NAND2_X1 _330_ (
  .A1(_068_),
  .A2(_070_),
  .ZN(_071_)
);

NAND3_X1 _331_ (
  .A1(_064_),
  .A2(_157_),
  .A3(_071_),
  .ZN(_072_)
);

NAND2_X1 _332_ (
  .A1(_167_),
  .A2(\coef[26] ),
  .ZN(_073_)
);

NAND2_X1 _333_ (
  .A1(_072_),
  .A2(_073_),
  .ZN(_004_)
);

NAND3_X1 _334_ (
  .A1(_050_),
  .A2(_051_),
  .A3(_121_),
  .ZN(_074_)
);

NAND2_X1 _335_ (
  .A1(_016_),
  .A2(_123_),
  .ZN(_075_)
);

INV_X1 _336_ (
  .A(_075_),
  .ZN(_076_)
);

AOI21_X1 _337_ (
  .A(_140_),
  .B1(_074_),
  .B2(_076_),
  .ZN(_077_)
);

INV_X1 _338_ (
  .A(_187_),
  .ZN(_078_)
);

NAND2_X1 _339_ (
  .A1(_078_),
  .A2(_132_),
  .ZN(_079_)
);

NAND2_X1 _340_ (
  .A1(_115_),
  .A2(_187_),
  .ZN(_080_)
);

NAND3_X1 _341_ (
  .A1(_079_),
  .A2(_080_),
  .A3(_120_),
  .ZN(_081_)
);

NAND2_X1 _342_ (
  .A1(_081_),
  .A2(_024_),
  .ZN(_082_)
);

NAND2_X1 _343_ (
  .A1(_082_),
  .A2(_162_),
  .ZN(_083_)
);

AOI21_X1 _344_ (
  .A(_167_),
  .B1(_077_),
  .B2(_083_),
  .ZN(_084_)
);

NAND2_X1 _345_ (
  .A1(_079_),
  .A2(_080_),
  .ZN(_085_)
);

NAND2_X1 _346_ (
  .A1(_085_),
  .A2(_126_),
  .ZN(_086_)
);

NAND2_X1 _347_ (
  .A1(_015_),
  .A2(_086_),
  .ZN(_087_)
);

NAND2_X1 _348_ (
  .A1(_087_),
  .A2(_165_),
  .ZN(_088_)
);

NAND3_X1 _349_ (
  .A1(_037_),
  .A2(_126_),
  .A3(_038_),
  .ZN(_089_)
);

NAND3_X1 _350_ (
  .A1(_089_),
  .A2(_162_),
  .A3(_025_),
  .ZN(_090_)
);

NAND3_X1 _351_ (
  .A1(_088_),
  .A2(_090_),
  .A3(_140_),
  .ZN(_091_)
);

NAND2_X1 _352_ (
  .A1(_084_),
  .A2(_091_),
  .ZN(_092_)
);

NAND2_X1 _353_ (
  .A1(_167_),
  .A2(\coef[13] ),
  .ZN(_093_)
);

NAND2_X1 _354_ (
  .A1(_092_),
  .A2(_093_),
  .ZN(_005_)
);

NOR2_X1 _355_ (
  .A1(_157_),
  .A2(\coef[28] ),
  .ZN(_094_)
);

NAND3_X1 _356_ (
  .A1(_086_),
  .A2(_165_),
  .A3(_025_),
  .ZN(_095_)
);

AOI21_X1 _357_ (
  .A(_140_),
  .B1(_161_),
  .B2(_162_),
  .ZN(_096_)
);

AOI21_X1 _358_ (
  .A(_167_),
  .B1(_095_),
  .B2(_096_),
  .ZN(_097_)
);

NAND3_X1 _359_ (
  .A1(_081_),
  .A2(_162_),
  .A3(_016_),
  .ZN(_098_)
);

OR2_X1 _360_ (
  .A1(_168_),
  .A2(_124_),
  .ZN(_099_)
);

NAND3_X1 _361_ (
  .A1(_098_),
  .A2(_140_),
  .A3(_099_),
  .ZN(_100_)
);

AOI21_X1 _362_ (
  .A(_094_),
  .B1(_097_),
  .B2(_100_),
  .ZN(_006_)
);

AOI21_X1 _363_ (
  .A(_140_),
  .B1(_086_),
  .B2(_154_),
  .ZN(_101_)
);

NAND2_X1 _364_ (
  .A1(_015_),
  .A2(_031_),
  .ZN(_102_)
);

NAND2_X1 _365_ (
  .A1(_102_),
  .A2(_165_),
  .ZN(_103_)
);

NAND2_X1 _366_ (
  .A1(_101_),
  .A2(_103_),
  .ZN(_104_)
);

AOI21_X1 _367_ (
  .A(_139_),
  .B1(_081_),
  .B2(_127_),
  .ZN(_105_)
);

NAND2_X1 _368_ (
  .A1(_044_),
  .A2(_024_),
  .ZN(_106_)
);

NAND2_X1 _369_ (
  .A1(_106_),
  .A2(_162_),
  .ZN(_107_)
);

NAND2_X1 _370_ (
  .A1(_105_),
  .A2(_107_),
  .ZN(_108_)
);

NAND3_X1 _371_ (
  .A1(_104_),
  .A2(_108_),
  .A3(_157_),
  .ZN(_109_)
);

NAND2_X1 _372_ (
  .A1(_167_),
  .A2(\coef[29] ),
  .ZN(_110_)
);

NAND2_X1 _373_ (
  .A1(_109_),
  .A2(_110_),
  .ZN(_007_)
);

NOR2_X1 _374_ (
  .A1(_157_),
  .A2(\coef[30] ),
  .ZN(_111_)
);

NOR2_X1 _375_ (
  .A1(_033_),
  .A2(_139_),
  .ZN(_112_)
);

NOR2_X1 _376_ (
  .A1(_112_),
  .A2(_046_),
  .ZN(_113_)
);

XNOR2_X1 _377_ (
  .A(_113_),
  .B(x[0]),
  .ZN(_114_)
);

AOI21_X1 _378_ (
  .A(_111_),
  .B1(_114_),
  .B2(_157_),
  .ZN(_008_)
);

HA_X1 _379_ (
  .A(_184_),
  .B(_185_),
  .CO(_186_),
  .S(_187_)
);

HA_X1 _380_ (
  .A(_184_),
  .B(_185_),
  .CO(_188_),
  .S(_189_)
);

HA_X1 _381_ (
  .A(_184_),
  .B(x[1]),
  .CO(_190_),
  .S(_191_)
);

HA_X1 _382_ (
  .A(_184_),
  .B(x[1]),
  .CO(_192_),
  .S(_193_)
);

HA_X1 _383_ (
  .A(x[0]),
  .B(_185_),
  .CO(_194_),
  .S(_195_)
);

HA_X1 _384_ (
  .A(x[0]),
  .B(_185_),
  .CO(_196_),
  .S(_197_)
);

HA_X1 _385_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_198_),
  .S(_199_)
);

HA_X1 _386_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_200_),
  .S(_201_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_183_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_182_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_181_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_180_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_179_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_178_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_177_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_176_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_175_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$785fe1ea8cdf428cbeb2f89081ee68c33feb7da2\dctu

module \$paramod$7911a3968b23dded19efefb86cf26bb44e3a7781\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _105_ (
  .A(x[1]),
  .ZN(_029_)
);

INV_X2 _106_ (
  .A(x[2]),
  .ZN(_030_)
);

NAND2_X4 _107_ (
  .A1(_029_),
  .A2(_030_),
  .ZN(_031_)
);

NAND2_X2 _108_ (
  .A1(x[1]),
  .A2(x[2]),
  .ZN(_032_)
);

NAND2_X2 _109_ (
  .A1(_031_),
  .A2(_032_),
  .ZN(_033_)
);

BUF_X4 _110_ (
  .A(y[0]),
  .Z(_034_)
);

INV_X2 _111_ (
  .A(_034_),
  .ZN(_035_)
);

NAND2_X2 _112_ (
  .A1(_033_),
  .A2(_035_),
  .ZN(_036_)
);

INV_X1 _113_ (
  .A(x[0]),
  .ZN(_037_)
);

NAND2_X1 _114_ (
  .A1(_030_),
  .A2(_037_),
  .ZN(_038_)
);

NAND2_X1 _115_ (
  .A1(x[2]),
  .A2(x[0]),
  .ZN(_039_)
);

NAND3_X2 _116_ (
  .A1(_038_),
  .A2(_034_),
  .A3(_039_),
  .ZN(_040_)
);

BUF_X4 _117_ (
  .A(y[1]),
  .Z(_041_)
);

NAND3_X1 _118_ (
  .A1(_036_),
  .A2(_040_),
  .A3(_041_),
  .ZN(_042_)
);

NAND3_X1 _119_ (
  .A1(_031_),
  .A2(_035_),
  .A3(_032_),
  .ZN(_043_)
);

INV_X2 _120_ (
  .A(_041_),
  .ZN(_044_)
);

NAND3_X1 _121_ (
  .A1(_043_),
  .A2(_040_),
  .A3(_044_),
  .ZN(_045_)
);

BUF_X4 _122_ (
  .A(y[2]),
  .Z(_046_)
);

NAND3_X1 _123_ (
  .A1(_042_),
  .A2(_045_),
  .A3(_046_),
  .ZN(_047_)
);

NAND2_X1 _124_ (
  .A1(_037_),
  .A2(x[2]),
  .ZN(_048_)
);

NAND2_X2 _125_ (
  .A1(_030_),
  .A2(x[0]),
  .ZN(_049_)
);

NAND2_X2 _126_ (
  .A1(_048_),
  .A2(_049_),
  .ZN(_050_)
);

NAND2_X4 _127_ (
  .A1(_050_),
  .A2(_035_),
  .ZN(_051_)
);

NAND3_X4 _128_ (
  .A1(_031_),
  .A2(_034_),
  .A3(_032_),
  .ZN(_052_)
);

NAND2_X4 _129_ (
  .A1(_051_),
  .A2(_052_),
  .ZN(_053_)
);

NAND2_X2 _130_ (
  .A1(_053_),
  .A2(_041_),
  .ZN(_054_)
);

NAND3_X2 _131_ (
  .A1(_048_),
  .A2(_049_),
  .A3(_035_),
  .ZN(_055_)
);

NAND3_X1 _132_ (
  .A1(_055_),
  .A2(_052_),
  .A3(_044_),
  .ZN(_056_)
);

INV_X2 _133_ (
  .A(_046_),
  .ZN(_057_)
);

NAND3_X1 _134_ (
  .A1(_054_),
  .A2(_056_),
  .A3(_057_),
  .ZN(_058_)
);

BUF_X1 _135_ (
  .A(ena),
  .Z(_059_)
);

BUF_X2 _136_ (
  .A(_059_),
  .Z(_060_)
);

NAND3_X1 _137_ (
  .A1(_047_),
  .A2(_058_),
  .A3(_060_),
  .ZN(_061_)
);

INV_X1 _138_ (
  .A(_059_),
  .ZN(_062_)
);

NAND2_X1 _139_ (
  .A1(_062_),
  .A2(\coef[21] ),
  .ZN(_063_)
);

NAND2_X1 _140_ (
  .A1(_061_),
  .A2(_063_),
  .ZN(_000_)
);

NAND3_X1 _141_ (
  .A1(_036_),
  .A2(_052_),
  .A3(_041_),
  .ZN(_064_)
);

INV_X1 _142_ (
  .A(_033_),
  .ZN(_065_)
);

AOI21_X1 _143_ (
  .A(_057_),
  .B1(_065_),
  .B2(_044_),
  .ZN(_066_)
);

NAND2_X1 _144_ (
  .A1(_064_),
  .A2(_066_),
  .ZN(_067_)
);

NAND3_X1 _145_ (
  .A1(_036_),
  .A2(_052_),
  .A3(_044_),
  .ZN(_068_)
);

AOI21_X1 _146_ (
  .A(_046_),
  .B1(_033_),
  .B2(_041_),
  .ZN(_069_)
);

NAND2_X1 _147_ (
  .A1(_068_),
  .A2(_069_),
  .ZN(_070_)
);

NAND3_X1 _148_ (
  .A1(_067_),
  .A2(_070_),
  .A3(_059_),
  .ZN(_071_)
);

INV_X1 _149_ (
  .A(\coef[22] ),
  .ZN(_072_)
);

OAI21_X1 _150_ (
  .A(_071_),
  .B1(_060_),
  .B2(_072_),
  .ZN(_001_)
);

NAND3_X1 _151_ (
  .A1(_043_),
  .A2(_040_),
  .A3(_041_),
  .ZN(_073_)
);

NAND3_X1 _152_ (
  .A1(_055_),
  .A2(_040_),
  .A3(_044_),
  .ZN(_074_)
);

NAND3_X1 _153_ (
  .A1(_073_),
  .A2(_074_),
  .A3(_046_),
  .ZN(_075_)
);

NAND2_X2 _154_ (
  .A1(_053_),
  .A2(_044_),
  .ZN(_076_)
);

NAND3_X1 _155_ (
  .A1(_055_),
  .A2(_040_),
  .A3(_041_),
  .ZN(_077_)
);

NAND3_X1 _156_ (
  .A1(_076_),
  .A2(_077_),
  .A3(_057_),
  .ZN(_078_)
);

NAND2_X1 _157_ (
  .A1(_075_),
  .A2(_078_),
  .ZN(_079_)
);

NAND2_X1 _158_ (
  .A1(_079_),
  .A2(_060_),
  .ZN(_080_)
);

NAND2_X1 _159_ (
  .A1(_062_),
  .A2(\coef[23] ),
  .ZN(_081_)
);

NAND2_X1 _160_ (
  .A1(_080_),
  .A2(_081_),
  .ZN(_002_)
);

NOR2_X1 _161_ (
  .A1(_059_),
  .A2(\coef[24] ),
  .ZN(_082_)
);

XNOR2_X1 _162_ (
  .A(_033_),
  .B(_041_),
  .ZN(_083_)
);

AOI21_X1 _163_ (
  .A(_082_),
  .B1(_083_),
  .B2(_060_),
  .ZN(_003_)
);

NAND3_X1 _164_ (
  .A1(_051_),
  .A2(_052_),
  .A3(_044_),
  .ZN(_084_)
);

NAND3_X1 _165_ (
  .A1(_077_),
  .A2(_084_),
  .A3(_046_),
  .ZN(_085_)
);

NAND2_X1 _166_ (
  .A1(_043_),
  .A2(_040_),
  .ZN(_086_)
);

NAND2_X1 _167_ (
  .A1(_086_),
  .A2(_041_),
  .ZN(_087_)
);

NAND3_X1 _168_ (
  .A1(_087_),
  .A2(_074_),
  .A3(_057_),
  .ZN(_088_)
);

NAND3_X1 _169_ (
  .A1(_085_),
  .A2(_088_),
  .A3(_060_),
  .ZN(_089_)
);

NAND2_X1 _170_ (
  .A1(_062_),
  .A2(\coef[25] ),
  .ZN(_090_)
);

NAND2_X1 _171_ (
  .A1(_089_),
  .A2(_090_),
  .ZN(_004_)
);

NAND2_X1 _172_ (
  .A1(_054_),
  .A2(_066_),
  .ZN(_091_)
);

NAND2_X1 _173_ (
  .A1(_045_),
  .A2(_069_),
  .ZN(_092_)
);

NAND3_X1 _174_ (
  .A1(_091_),
  .A2(_092_),
  .A3(_059_),
  .ZN(_093_)
);

INV_X1 _175_ (
  .A(\coef[26] ),
  .ZN(_094_)
);

OAI21_X1 _176_ (
  .A(_093_),
  .B1(_060_),
  .B2(_094_),
  .ZN(_005_)
);

NAND3_X1 _177_ (
  .A1(_055_),
  .A2(_052_),
  .A3(_041_),
  .ZN(_010_)
);

NAND3_X1 _178_ (
  .A1(_076_),
  .A2(_010_),
  .A3(_046_),
  .ZN(_011_)
);

NAND3_X1 _179_ (
  .A1(_036_),
  .A2(_040_),
  .A3(_044_),
  .ZN(_012_)
);

NAND3_X1 _180_ (
  .A1(_073_),
  .A2(_012_),
  .A3(_057_),
  .ZN(_013_)
);

NAND2_X1 _181_ (
  .A1(_011_),
  .A2(_013_),
  .ZN(_014_)
);

NAND2_X1 _182_ (
  .A1(_014_),
  .A2(_060_),
  .ZN(_015_)
);

NAND2_X1 _183_ (
  .A1(_062_),
  .A2(\coef[27] ),
  .ZN(_016_)
);

NAND2_X1 _184_ (
  .A1(_015_),
  .A2(_016_),
  .ZN(_006_)
);

NOR2_X1 _185_ (
  .A1(_059_),
  .A2(\coef[28] ),
  .ZN(_017_)
);

OAI21_X1 _186_ (
  .A(_044_),
  .B1(_035_),
  .B2(_057_),
  .ZN(_018_)
);

OAI21_X1 _187_ (
  .A(_018_),
  .B1(_034_),
  .B2(_046_),
  .ZN(_019_)
);

XOR2_X1 _188_ (
  .A(_019_),
  .B(_050_),
  .Z(_020_)
);

AOI21_X1 _189_ (
  .A(_017_),
  .B1(_020_),
  .B2(_060_),
  .ZN(_007_)
);

NAND3_X1 _190_ (
  .A1(_045_),
  .A2(_064_),
  .A3(_046_),
  .ZN(_021_)
);

NAND3_X1 _191_ (
  .A1(_054_),
  .A2(_068_),
  .A3(_057_),
  .ZN(_022_)
);

NAND3_X1 _192_ (
  .A1(_021_),
  .A2(_022_),
  .A3(_060_),
  .ZN(_023_)
);

NAND2_X1 _193_ (
  .A1(_062_),
  .A2(\coef[15] ),
  .ZN(_024_)
);

NAND2_X1 _194_ (
  .A1(_023_),
  .A2(_024_),
  .ZN(_008_)
);

NOR2_X1 _195_ (
  .A1(_059_),
  .A2(\coef[30] ),
  .ZN(_025_)
);

OAI21_X1 _196_ (
  .A(_044_),
  .B1(_034_),
  .B2(_046_),
  .ZN(_026_)
);

OAI21_X1 _197_ (
  .A(_026_),
  .B1(_035_),
  .B2(_057_),
  .ZN(_027_)
);

XNOR2_X1 _198_ (
  .A(_027_),
  .B(_050_),
  .ZN(_028_)
);

AOI21_X1 _199_ (
  .A(_025_),
  .B1(_028_),
  .B2(_060_),
  .ZN(_009_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_104_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_103_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_102_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_101_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_100_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_099_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_098_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_097_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_096_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_095_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$7911a3968b23dded19efefb86cf26bb44e3a7781\dctu

module \$paramod$826cb5d104d530340b1f58495d2410742b2c32fe\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _189_ (
  .A(x[0]),
  .ZN(_171_)
);

INV_X1 _190_ (
  .A(x[1]),
  .ZN(_172_)
);

BUF_X1 _191_ (
  .A(ena),
  .Z(_103_)
);

NOR2_X1 _192_ (
  .A1(\coef[21] ),
  .A2(_103_),
  .ZN(_104_)
);

BUF_X8 _193_ (
  .A(x[2]),
  .Z(_105_)
);

INV_X8 _194_ (
  .A(_105_),
  .ZN(_106_)
);

INV_X1 _195_ (
  .A(_185_),
  .ZN(_107_)
);

NAND2_X2 _196_ (
  .A1(_106_),
  .A2(_107_),
  .ZN(_108_)
);

BUF_X16 _197_ (
  .A(_105_),
  .Z(_109_)
);

NAND2_X4 _198_ (
  .A1(_109_),
  .A2(_175_),
  .ZN(_110_)
);

NAND2_X4 _199_ (
  .A1(_108_),
  .A2(_110_),
  .ZN(_111_)
);

BUF_X4 _200_ (
  .A(y[0]),
  .Z(_112_)
);

INV_X8 _201_ (
  .A(_112_),
  .ZN(_113_)
);

NAND2_X4 _202_ (
  .A1(_111_),
  .A2(_113_),
  .ZN(_114_)
);

NAND2_X1 _203_ (
  .A1(_106_),
  .A2(_181_),
  .ZN(_115_)
);

INV_X1 _204_ (
  .A(_179_),
  .ZN(_116_)
);

NAND2_X1 _205_ (
  .A1(_116_),
  .A2(_109_),
  .ZN(_117_)
);

BUF_X4 _206_ (
  .A(_112_),
  .Z(_118_)
);

NAND3_X1 _207_ (
  .A1(_115_),
  .A2(_117_),
  .A3(_118_),
  .ZN(_119_)
);

NAND2_X1 _208_ (
  .A1(_114_),
  .A2(_119_),
  .ZN(_120_)
);

BUF_X4 _209_ (
  .A(y[2]),
  .Z(_121_)
);

INV_X2 _210_ (
  .A(_121_),
  .ZN(_122_)
);

BUF_X4 _211_ (
  .A(y[1]),
  .Z(_123_)
);

NOR2_X4 _212_ (
  .A1(_122_),
  .A2(_123_),
  .ZN(_124_)
);

NAND2_X1 _213_ (
  .A1(_120_),
  .A2(_124_),
  .ZN(_125_)
);

INV_X1 _214_ (
  .A(_181_),
  .ZN(_126_)
);

NAND2_X2 _215_ (
  .A1(_106_),
  .A2(_126_),
  .ZN(_127_)
);

BUF_X4 _216_ (
  .A(_113_),
  .Z(_128_)
);

NAND2_X4 _217_ (
  .A1(_109_),
  .A2(_179_),
  .ZN(_129_)
);

NAND3_X1 _218_ (
  .A1(_127_),
  .A2(_128_),
  .A3(_129_),
  .ZN(_130_)
);

NAND3_X2 _219_ (
  .A1(_108_),
  .A2(_118_),
  .A3(_110_),
  .ZN(_131_)
);

INV_X2 _220_ (
  .A(_123_),
  .ZN(_132_)
);

NOR2_X4 _221_ (
  .A1(_132_),
  .A2(_121_),
  .ZN(_133_)
);

NAND3_X1 _222_ (
  .A1(_130_),
  .A2(_131_),
  .A3(_133_),
  .ZN(_134_)
);

NAND2_X1 _223_ (
  .A1(_125_),
  .A2(_134_),
  .ZN(_135_)
);

NOR2_X2 _224_ (
  .A1(_123_),
  .A2(_121_),
  .ZN(_136_)
);

INV_X1 _225_ (
  .A(_136_),
  .ZN(_137_)
);

OR2_X4 _226_ (
  .A1(_187_),
  .A2(_105_),
  .ZN(_138_)
);

NAND2_X1 _227_ (
  .A1(_105_),
  .A2(_173_),
  .ZN(_139_)
);

NAND3_X1 _228_ (
  .A1(_138_),
  .A2(_128_),
  .A3(_139_),
  .ZN(_140_)
);

INV_X1 _229_ (
  .A(_183_),
  .ZN(_141_)
);

NAND2_X2 _230_ (
  .A1(_106_),
  .A2(_141_),
  .ZN(_142_)
);

NAND2_X4 _231_ (
  .A1(_109_),
  .A2(_177_),
  .ZN(_143_)
);

NAND3_X2 _232_ (
  .A1(_142_),
  .A2(_118_),
  .A3(_143_),
  .ZN(_144_)
);

AOI21_X1 _233_ (
  .A(_137_),
  .B1(_140_),
  .B2(_144_),
  .ZN(_145_)
);

NOR2_X2 _234_ (
  .A1(_135_),
  .A2(_145_),
  .ZN(_146_)
);

NAND2_X1 _235_ (
  .A1(_123_),
  .A2(_121_),
  .ZN(_147_)
);

NAND3_X1 _236_ (
  .A1(_138_),
  .A2(_118_),
  .A3(_139_),
  .ZN(_148_)
);

NAND3_X1 _237_ (
  .A1(_142_),
  .A2(_128_),
  .A3(_143_),
  .ZN(_149_)
);

AOI21_X1 _238_ (
  .A(_147_),
  .B1(_148_),
  .B2(_149_),
  .ZN(_150_)
);

INV_X1 _239_ (
  .A(_103_),
  .ZN(_151_)
);

NOR2_X1 _240_ (
  .A1(_150_),
  .A2(_151_),
  .ZN(_152_)
);

AOI21_X2 _241_ (
  .A(_104_),
  .B1(_146_),
  .B2(_152_),
  .ZN(_000_)
);

BUF_X4 _242_ (
  .A(_103_),
  .Z(_153_)
);

XNOR2_X1 _243_ (
  .A(_112_),
  .B(_121_),
  .ZN(_154_)
);

NAND2_X2 _244_ (
  .A1(_109_),
  .A2(_187_),
  .ZN(_155_)
);

INV_X1 _245_ (
  .A(_173_),
  .ZN(_156_)
);

NAND2_X1 _246_ (
  .A1(_106_),
  .A2(_156_),
  .ZN(_157_)
);

AOI21_X1 _247_ (
  .A(_154_),
  .B1(_155_),
  .B2(_157_),
  .ZN(_158_)
);

INV_X1 _248_ (
  .A(_175_),
  .ZN(_159_)
);

NAND2_X1 _249_ (
  .A1(_106_),
  .A2(_159_),
  .ZN(_160_)
);

NAND2_X2 _250_ (
  .A1(_109_),
  .A2(_185_),
  .ZN(_010_)
);

NAND2_X2 _251_ (
  .A1(_160_),
  .A2(_010_),
  .ZN(_011_)
);

INV_X1 _252_ (
  .A(_011_),
  .ZN(_012_)
);

AND2_X1 _253_ (
  .A1(_012_),
  .A2(_154_),
  .ZN(_013_)
);

OAI21_X1 _254_ (
  .A(_153_),
  .B1(_158_),
  .B2(_013_),
  .ZN(_014_)
);

INV_X1 _255_ (
  .A(\coef[22] ),
  .ZN(_015_)
);

OAI21_X1 _256_ (
  .A(_014_),
  .B1(_153_),
  .B2(_015_),
  .ZN(_001_)
);

NAND2_X2 _257_ (
  .A1(_138_),
  .A2(_139_),
  .ZN(_016_)
);

NAND2_X1 _258_ (
  .A1(_016_),
  .A2(_113_),
  .ZN(_017_)
);

OAI21_X1 _259_ (
  .A(_123_),
  .B1(_113_),
  .B2(x[0]),
  .ZN(_018_)
);

INV_X1 _260_ (
  .A(_018_),
  .ZN(_019_)
);

NAND2_X1 _261_ (
  .A1(_017_),
  .A2(_019_),
  .ZN(_020_)
);

AOI21_X1 _262_ (
  .A(_123_),
  .B1(_113_),
  .B2(x[0]),
  .ZN(_021_)
);

NAND2_X1 _263_ (
  .A1(_131_),
  .A2(_021_),
  .ZN(_022_)
);

NAND2_X1 _264_ (
  .A1(_020_),
  .A2(_022_),
  .ZN(_023_)
);

NAND2_X1 _265_ (
  .A1(_023_),
  .A2(_122_),
  .ZN(_024_)
);

NAND2_X1 _266_ (
  .A1(_148_),
  .A2(_021_),
  .ZN(_025_)
);

NAND2_X2 _267_ (
  .A1(_114_),
  .A2(_019_),
  .ZN(_026_)
);

NAND3_X1 _268_ (
  .A1(_025_),
  .A2(_026_),
  .A3(_121_),
  .ZN(_027_)
);

NAND2_X1 _269_ (
  .A1(_024_),
  .A2(_027_),
  .ZN(_028_)
);

NAND2_X2 _270_ (
  .A1(_028_),
  .A2(_153_),
  .ZN(_029_)
);

NAND2_X1 _271_ (
  .A1(_151_),
  .A2(\coef[23] ),
  .ZN(_030_)
);

NAND2_X2 _272_ (
  .A1(_029_),
  .A2(_030_),
  .ZN(_002_)
);

NOR2_X1 _273_ (
  .A1(_153_),
  .A2(\coef[24] ),
  .ZN(_031_)
);

XNOR2_X1 _274_ (
  .A(_154_),
  .B(_172_),
  .ZN(_032_)
);

AOI21_X1 _275_ (
  .A(_031_),
  .B1(_032_),
  .B2(_153_),
  .ZN(_003_)
);

NOR2_X1 _276_ (
  .A1(_103_),
  .A2(\coef[25] ),
  .ZN(_033_)
);

NAND2_X4 _277_ (
  .A1(_142_),
  .A2(_143_),
  .ZN(_034_)
);

NAND2_X1 _278_ (
  .A1(_034_),
  .A2(_118_),
  .ZN(_035_)
);

INV_X1 _279_ (
  .A(_174_),
  .ZN(_036_)
);

NAND2_X2 _280_ (
  .A1(_106_),
  .A2(_036_),
  .ZN(_037_)
);

NAND2_X4 _281_ (
  .A1(_109_),
  .A2(_174_),
  .ZN(_038_)
);

NAND2_X4 _282_ (
  .A1(_037_),
  .A2(_038_),
  .ZN(_039_)
);

NAND2_X4 _283_ (
  .A1(_039_),
  .A2(_113_),
  .ZN(_040_)
);

NAND3_X1 _284_ (
  .A1(_035_),
  .A2(_040_),
  .A3(_136_),
  .ZN(_041_)
);

NAND3_X4 _285_ (
  .A1(_037_),
  .A2(_118_),
  .A3(_038_),
  .ZN(_042_)
);

NAND3_X1 _286_ (
  .A1(_130_),
  .A2(_042_),
  .A3(_133_),
  .ZN(_043_)
);

NAND2_X1 _287_ (
  .A1(_041_),
  .A2(_043_),
  .ZN(_044_)
);

AOI21_X1 _288_ (
  .A(_147_),
  .B1(_149_),
  .B2(_042_),
  .ZN(_045_)
);

NOR2_X2 _289_ (
  .A1(_044_),
  .A2(_045_),
  .ZN(_046_)
);

NAND2_X1 _290_ (
  .A1(_040_),
  .A2(_119_),
  .ZN(_047_)
);

AOI21_X1 _291_ (
  .A(_151_),
  .B1(_047_),
  .B2(_124_),
  .ZN(_048_)
);

AOI21_X2 _292_ (
  .A(_033_),
  .B1(_046_),
  .B2(_048_),
  .ZN(_004_)
);

NOR2_X1 _293_ (
  .A1(_153_),
  .A2(\coef[26] ),
  .ZN(_049_)
);

OAI21_X1 _294_ (
  .A(_123_),
  .B1(_109_),
  .B2(_112_),
  .ZN(_050_)
);

INV_X1 _295_ (
  .A(_050_),
  .ZN(_051_)
);

AOI21_X1 _296_ (
  .A(_122_),
  .B1(_144_),
  .B2(_051_),
  .ZN(_052_)
);

NAND2_X2 _297_ (
  .A1(_127_),
  .A2(_129_),
  .ZN(_053_)
);

NAND2_X1 _298_ (
  .A1(_053_),
  .A2(_128_),
  .ZN(_054_)
);

OAI21_X1 _299_ (
  .A(_132_),
  .B1(_106_),
  .B2(_113_),
  .ZN(_055_)
);

INV_X1 _300_ (
  .A(_055_),
  .ZN(_056_)
);

NAND2_X1 _301_ (
  .A1(_054_),
  .A2(_056_),
  .ZN(_057_)
);

AOI21_X1 _302_ (
  .A(_151_),
  .B1(_052_),
  .B2(_057_),
  .ZN(_058_)
);

NAND3_X2 _303_ (
  .A1(_127_),
  .A2(_118_),
  .A3(_129_),
  .ZN(_059_)
);

NAND2_X1 _304_ (
  .A1(_059_),
  .A2(_051_),
  .ZN(_060_)
);

NAND2_X2 _305_ (
  .A1(_034_),
  .A2(_128_),
  .ZN(_061_)
);

INV_X1 _306_ (
  .A(_061_),
  .ZN(_062_)
);

OAI21_X2 _307_ (
  .A(_060_),
  .B1(_062_),
  .B2(_055_),
  .ZN(_063_)
);

NAND2_X1 _308_ (
  .A1(_063_),
  .A2(_122_),
  .ZN(_064_)
);

AOI21_X2 _309_ (
  .A(_049_),
  .B1(_058_),
  .B2(_064_),
  .ZN(_005_)
);

NOR2_X1 _310_ (
  .A1(_153_),
  .A2(\coef[27] ),
  .ZN(_065_)
);

INV_X1 _311_ (
  .A(_177_),
  .ZN(_066_)
);

NAND2_X1 _312_ (
  .A1(_106_),
  .A2(_066_),
  .ZN(_067_)
);

NAND2_X1 _313_ (
  .A1(_109_),
  .A2(_183_),
  .ZN(_068_)
);

NAND3_X1 _314_ (
  .A1(_067_),
  .A2(_118_),
  .A3(_068_),
  .ZN(_069_)
);

NAND3_X1 _315_ (
  .A1(_157_),
  .A2(_128_),
  .A3(_155_),
  .ZN(_070_)
);

NAND3_X1 _316_ (
  .A1(_069_),
  .A2(_070_),
  .A3(_133_),
  .ZN(_071_)
);

NAND3_X1 _317_ (
  .A1(_067_),
  .A2(_128_),
  .A3(_068_),
  .ZN(_072_)
);

NAND3_X1 _318_ (
  .A1(_157_),
  .A2(_118_),
  .A3(_155_),
  .ZN(_073_)
);

NAND3_X1 _319_ (
  .A1(_072_),
  .A2(_073_),
  .A3(_124_),
  .ZN(_074_)
);

NAND2_X1 _320_ (
  .A1(_071_),
  .A2(_074_),
  .ZN(_075_)
);

NAND2_X1 _321_ (
  .A1(_012_),
  .A2(_128_),
  .ZN(_076_)
);

NAND2_X1 _322_ (
  .A1(_106_),
  .A2(_116_),
  .ZN(_077_)
);

NAND2_X1 _323_ (
  .A1(_109_),
  .A2(_181_),
  .ZN(_078_)
);

NAND3_X1 _324_ (
  .A1(_077_),
  .A2(_118_),
  .A3(_078_),
  .ZN(_079_)
);

AOI21_X1 _325_ (
  .A(_147_),
  .B1(_076_),
  .B2(_079_),
  .ZN(_080_)
);

NOR2_X1 _326_ (
  .A1(_075_),
  .A2(_080_),
  .ZN(_081_)
);

NAND3_X1 _327_ (
  .A1(_077_),
  .A2(_128_),
  .A3(_078_),
  .ZN(_082_)
);

OAI21_X1 _328_ (
  .A(_082_),
  .B1(_128_),
  .B2(_011_),
  .ZN(_083_)
);

AOI21_X1 _329_ (
  .A(_151_),
  .B1(_083_),
  .B2(_136_),
  .ZN(_084_)
);

AOI21_X2 _330_ (
  .A(_065_),
  .B1(_081_),
  .B2(_084_),
  .ZN(_006_)
);

NOR2_X2 _331_ (
  .A1(_133_),
  .A2(_124_),
  .ZN(_085_)
);

AOI21_X1 _332_ (
  .A(_151_),
  .B1(_085_),
  .B2(_016_),
  .ZN(_086_)
);

OAI21_X1 _333_ (
  .A(_086_),
  .B1(_111_),
  .B2(_085_),
  .ZN(_087_)
);

INV_X1 _334_ (
  .A(\coef[28] ),
  .ZN(_088_)
);

OAI21_X1 _335_ (
  .A(_087_),
  .B1(_153_),
  .B2(_088_),
  .ZN(_007_)
);

NOR2_X1 _336_ (
  .A1(_153_),
  .A2(\coef[15] ),
  .ZN(_089_)
);

NAND2_X2 _337_ (
  .A1(_040_),
  .A2(_144_),
  .ZN(_090_)
);

NAND2_X2 _338_ (
  .A1(_090_),
  .A2(_136_),
  .ZN(_091_)
);

NAND2_X2 _339_ (
  .A1(_091_),
  .A2(_103_),
  .ZN(_092_)
);

INV_X1 _340_ (
  .A(_133_),
  .ZN(_093_)
);

AOI21_X1 _341_ (
  .A(_093_),
  .B1(_054_),
  .B2(_042_),
  .ZN(_094_)
);

NOR2_X2 _342_ (
  .A1(_092_),
  .A2(_094_),
  .ZN(_095_)
);

NAND3_X1 _343_ (
  .A1(_061_),
  .A2(_042_),
  .A3(_123_),
  .ZN(_096_)
);

NAND3_X2 _344_ (
  .A1(_040_),
  .A2(_059_),
  .A3(_132_),
  .ZN(_097_)
);

NAND2_X1 _345_ (
  .A1(_096_),
  .A2(_097_),
  .ZN(_098_)
);

NAND2_X1 _346_ (
  .A1(_098_),
  .A2(_121_),
  .ZN(_099_)
);

AOI21_X2 _347_ (
  .A(_089_),
  .B1(_095_),
  .B2(_099_),
  .ZN(_008_)
);

AOI21_X1 _348_ (
  .A(_151_),
  .B1(_085_),
  .B2(_034_),
  .ZN(_100_)
);

OAI21_X1 _349_ (
  .A(_100_),
  .B1(_053_),
  .B2(_085_),
  .ZN(_101_)
);

INV_X1 _350_ (
  .A(\coef[30] ),
  .ZN(_102_)
);

OAI21_X1 _351_ (
  .A(_101_),
  .B1(_153_),
  .B2(_102_),
  .ZN(_009_)
);

HA_X1 _352_ (
  .A(_171_),
  .B(_172_),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _353_ (
  .A(_171_),
  .B(_172_),
  .CO(_175_),
  .S(_176_)
);

HA_X1 _354_ (
  .A(_171_),
  .B(x[1]),
  .CO(_177_),
  .S(_178_)
);

HA_X1 _355_ (
  .A(_171_),
  .B(x[1]),
  .CO(_179_),
  .S(_180_)
);

HA_X1 _356_ (
  .A(x[0]),
  .B(_172_),
  .CO(_181_),
  .S(_182_)
);

HA_X1 _357_ (
  .A(x[0]),
  .B(_172_),
  .CO(_183_),
  .S(_184_)
);

HA_X1 _358_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_185_),
  .S(_186_)
);

HA_X1 _359_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_187_),
  .S(_188_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_170_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_169_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_168_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_167_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_166_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_165_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_164_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_163_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_162_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_161_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$826cb5d104d530340b1f58495d2410742b2c32fe\dctu

module \$paramod$0c5a5bd6be4ed818deaac08b02afbddb6897ffee\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

BUF_X2 _178_ (
  .A(x[0]),
  .Z(_093_)
);

INV_X1 _179_ (
  .A(_093_),
  .ZN(_160_)
);

INV_X1 _180_ (
  .A(x[1]),
  .ZN(_161_)
);

INV_X2 _181_ (
  .A(x[2]),
  .ZN(_094_)
);

NAND2_X1 _182_ (
  .A1(_094_),
  .A2(_163_),
  .ZN(_095_)
);

INV_X1 _183_ (
  .A(_163_),
  .ZN(_096_)
);

BUF_X4 _184_ (
  .A(x[2]),
  .Z(_097_)
);

NAND2_X1 _185_ (
  .A1(_096_),
  .A2(_097_),
  .ZN(_098_)
);

BUF_X4 _186_ (
  .A(y[0]),
  .Z(_099_)
);

INV_X8 _187_ (
  .A(_099_),
  .ZN(_100_)
);

NAND3_X1 _188_ (
  .A1(_095_),
  .A2(_098_),
  .A3(_100_),
  .ZN(_101_)
);

NOR2_X2 _189_ (
  .A1(_100_),
  .A2(_093_),
  .ZN(_102_)
);

BUF_X4 _190_ (
  .A(y[1]),
  .Z(_103_)
);

NOR2_X1 _191_ (
  .A1(_102_),
  .A2(_103_),
  .ZN(_104_)
);

NAND2_X1 _192_ (
  .A1(_101_),
  .A2(_104_),
  .ZN(_105_)
);

BUF_X8 _193_ (
  .A(_094_),
  .Z(_106_)
);

NAND2_X2 _194_ (
  .A1(_106_),
  .A2(_096_),
  .ZN(_107_)
);

BUF_X8 _195_ (
  .A(_099_),
  .Z(_108_)
);

NAND2_X1 _196_ (
  .A1(_097_),
  .A2(_163_),
  .ZN(_109_)
);

NAND3_X2 _197_ (
  .A1(_107_),
  .A2(_108_),
  .A3(_109_),
  .ZN(_110_)
);

NAND2_X1 _198_ (
  .A1(_100_),
  .A2(_093_),
  .ZN(_111_)
);

NAND2_X1 _199_ (
  .A1(_111_),
  .A2(_103_),
  .ZN(_112_)
);

INV_X1 _200_ (
  .A(_112_),
  .ZN(_113_)
);

NAND2_X1 _201_ (
  .A1(_110_),
  .A2(_113_),
  .ZN(_114_)
);

NAND2_X1 _202_ (
  .A1(_105_),
  .A2(_114_),
  .ZN(_115_)
);

BUF_X4 _203_ (
  .A(y[2]),
  .Z(_116_)
);

NAND2_X1 _204_ (
  .A1(_115_),
  .A2(_116_),
  .ZN(_117_)
);

INV_X4 _205_ (
  .A(_116_),
  .ZN(_118_)
);

NAND3_X1 _206_ (
  .A1(_105_),
  .A2(_114_),
  .A3(_118_),
  .ZN(_119_)
);

BUF_X1 _207_ (
  .A(ena),
  .Z(_120_)
);

BUF_X2 _208_ (
  .A(_120_),
  .Z(_121_)
);

NAND3_X1 _209_ (
  .A1(_117_),
  .A2(_119_),
  .A3(_121_),
  .ZN(_122_)
);

INV_X1 _210_ (
  .A(_120_),
  .ZN(_123_)
);

NAND2_X1 _211_ (
  .A1(_123_),
  .A2(\coef[21] ),
  .ZN(_124_)
);

NAND2_X1 _212_ (
  .A1(_122_),
  .A2(_124_),
  .ZN(_000_)
);

NOR2_X1 _213_ (
  .A1(_120_),
  .A2(\coef[22] ),
  .ZN(_125_)
);

XNOR2_X2 _214_ (
  .A(_108_),
  .B(_116_),
  .ZN(_126_)
);

XNOR2_X1 _215_ (
  .A(_126_),
  .B(_106_),
  .ZN(_127_)
);

AOI21_X1 _216_ (
  .A(_125_),
  .B1(_127_),
  .B2(_121_),
  .ZN(_001_)
);

NOR2_X1 _217_ (
  .A1(_120_),
  .A2(\coef[23] ),
  .ZN(_128_)
);

INV_X1 _218_ (
  .A(_162_),
  .ZN(_129_)
);

NAND2_X1 _219_ (
  .A1(_094_),
  .A2(_129_),
  .ZN(_130_)
);

NAND2_X1 _220_ (
  .A1(x[2]),
  .A2(_176_),
  .ZN(_131_)
);

NAND2_X1 _221_ (
  .A1(_130_),
  .A2(_131_),
  .ZN(_132_)
);

NAND2_X1 _222_ (
  .A1(_132_),
  .A2(_100_),
  .ZN(_133_)
);

NAND2_X1 _223_ (
  .A1(_133_),
  .A2(_110_),
  .ZN(_134_)
);

NOR2_X4 _224_ (
  .A1(_118_),
  .A2(y[1]),
  .ZN(_135_)
);

NAND2_X1 _225_ (
  .A1(_134_),
  .A2(_135_),
  .ZN(_136_)
);

NAND2_X1 _226_ (
  .A1(_136_),
  .A2(_120_),
  .ZN(_137_)
);

NAND2_X1 _227_ (
  .A1(_103_),
  .A2(_116_),
  .ZN(_138_)
);

NAND2_X1 _228_ (
  .A1(_106_),
  .A2(_164_),
  .ZN(_139_)
);

INV_X1 _229_ (
  .A(_174_),
  .ZN(_140_)
);

NAND2_X1 _230_ (
  .A1(_140_),
  .A2(_097_),
  .ZN(_141_)
);

NAND2_X1 _231_ (
  .A1(_139_),
  .A2(_141_),
  .ZN(_142_)
);

NAND2_X1 _232_ (
  .A1(_142_),
  .A2(_108_),
  .ZN(_143_)
);

AOI21_X1 _233_ (
  .A(_138_),
  .B1(_143_),
  .B2(_101_),
  .ZN(_144_)
);

NOR2_X1 _234_ (
  .A1(_137_),
  .A2(_144_),
  .ZN(_145_)
);

NAND3_X1 _235_ (
  .A1(_130_),
  .A2(_108_),
  .A3(_131_),
  .ZN(_146_)
);

NAND3_X1 _236_ (
  .A1(_101_),
  .A2(_146_),
  .A3(_103_),
  .ZN(_147_)
);

NAND3_X1 _237_ (
  .A1(_139_),
  .A2(_141_),
  .A3(_100_),
  .ZN(_148_)
);

INV_X1 _238_ (
  .A(_103_),
  .ZN(_149_)
);

NAND3_X1 _239_ (
  .A1(_148_),
  .A2(_110_),
  .A3(_149_),
  .ZN(_010_)
);

NAND2_X1 _240_ (
  .A1(_147_),
  .A2(_010_),
  .ZN(_011_)
);

NAND2_X1 _241_ (
  .A1(_011_),
  .A2(_118_),
  .ZN(_012_)
);

AOI21_X2 _242_ (
  .A(_128_),
  .B1(_145_),
  .B2(_012_),
  .ZN(_002_)
);

NAND2_X1 _243_ (
  .A1(_123_),
  .A2(\coef[24] ),
  .ZN(_013_)
);

NAND2_X1 _244_ (
  .A1(_106_),
  .A2(_140_),
  .ZN(_014_)
);

NAND2_X1 _245_ (
  .A1(_097_),
  .A2(_164_),
  .ZN(_015_)
);

NAND3_X1 _246_ (
  .A1(_126_),
  .A2(_014_),
  .A3(_015_),
  .ZN(_016_)
);

NAND2_X1 _247_ (
  .A1(_016_),
  .A2(_121_),
  .ZN(_017_)
);

NAND2_X1 _248_ (
  .A1(_106_),
  .A2(_176_),
  .ZN(_018_)
);

OAI21_X1 _249_ (
  .A(_018_),
  .B1(_106_),
  .B2(_162_),
  .ZN(_019_)
);

NOR2_X1 _250_ (
  .A1(_019_),
  .A2(_126_),
  .ZN(_020_)
);

OAI21_X1 _251_ (
  .A(_013_),
  .B1(_017_),
  .B2(_020_),
  .ZN(_003_)
);

NAND2_X2 _252_ (
  .A1(_106_),
  .A2(_166_),
  .ZN(_021_)
);

INV_X1 _253_ (
  .A(_172_),
  .ZN(_022_)
);

NAND2_X1 _254_ (
  .A1(_022_),
  .A2(_097_),
  .ZN(_023_)
);

NAND3_X1 _255_ (
  .A1(_021_),
  .A2(_023_),
  .A3(_100_),
  .ZN(_024_)
);

NAND2_X1 _256_ (
  .A1(_093_),
  .A2(_108_),
  .ZN(_025_)
);

NAND2_X1 _257_ (
  .A1(_024_),
  .A2(_025_),
  .ZN(_026_)
);

NOR2_X1 _258_ (
  .A1(_103_),
  .A2(_116_),
  .ZN(_027_)
);

NAND2_X1 _259_ (
  .A1(_026_),
  .A2(_027_),
  .ZN(_028_)
);

NAND3_X1 _260_ (
  .A1(_021_),
  .A2(_023_),
  .A3(_108_),
  .ZN(_029_)
);

NAND2_X1 _261_ (
  .A1(_029_),
  .A2(_111_),
  .ZN(_030_)
);

INV_X1 _262_ (
  .A(_138_),
  .ZN(_031_)
);

NAND2_X1 _263_ (
  .A1(_030_),
  .A2(_031_),
  .ZN(_032_)
);

INV_X1 _264_ (
  .A(_168_),
  .ZN(_033_)
);

NAND2_X4 _265_ (
  .A1(_106_),
  .A2(_033_),
  .ZN(_034_)
);

NAND2_X2 _266_ (
  .A1(_097_),
  .A2(_170_),
  .ZN(_035_)
);

NAND3_X1 _267_ (
  .A1(_034_),
  .A2(_108_),
  .A3(_035_),
  .ZN(_036_)
);

NOR2_X1 _268_ (
  .A1(_093_),
  .A2(_099_),
  .ZN(_037_)
);

INV_X1 _269_ (
  .A(_037_),
  .ZN(_038_)
);

NAND2_X1 _270_ (
  .A1(_036_),
  .A2(_038_),
  .ZN(_039_)
);

NAND2_X1 _271_ (
  .A1(_118_),
  .A2(y[1]),
  .ZN(_040_)
);

INV_X1 _272_ (
  .A(_040_),
  .ZN(_041_)
);

NAND2_X1 _273_ (
  .A1(_039_),
  .A2(_041_),
  .ZN(_042_)
);

NAND3_X1 _274_ (
  .A1(_028_),
  .A2(_032_),
  .A3(_042_),
  .ZN(_043_)
);

NAND3_X2 _275_ (
  .A1(_034_),
  .A2(_100_),
  .A3(_035_),
  .ZN(_044_)
);

INV_X1 _276_ (
  .A(_102_),
  .ZN(_045_)
);

AND2_X1 _277_ (
  .A1(_044_),
  .A2(_045_),
  .ZN(_046_)
);

INV_X1 _278_ (
  .A(_135_),
  .ZN(_047_)
);

OAI21_X1 _279_ (
  .A(_120_),
  .B1(_046_),
  .B2(_047_),
  .ZN(_048_)
);

NOR2_X1 _280_ (
  .A1(_043_),
  .A2(_048_),
  .ZN(_049_)
);

NOR2_X1 _281_ (
  .A1(_121_),
  .A2(\coef[25] ),
  .ZN(_050_)
);

NOR2_X2 _282_ (
  .A1(_049_),
  .A2(_050_),
  .ZN(_004_)
);

NAND2_X1 _283_ (
  .A1(_123_),
  .A2(\coef[26] ),
  .ZN(_051_)
);

NAND2_X1 _284_ (
  .A1(_106_),
  .A2(_170_),
  .ZN(_052_)
);

NAND2_X1 _285_ (
  .A1(_033_),
  .A2(_097_),
  .ZN(_053_)
);

NAND3_X1 _286_ (
  .A1(_052_),
  .A2(_053_),
  .A3(_100_),
  .ZN(_054_)
);

NAND3_X1 _287_ (
  .A1(_054_),
  .A2(_103_),
  .A3(_025_),
  .ZN(_055_)
);

NOR2_X1 _288_ (
  .A1(_037_),
  .A2(_103_),
  .ZN(_056_)
);

NAND2_X1 _289_ (
  .A1(_097_),
  .A2(_166_),
  .ZN(_057_)
);

OAI21_X1 _290_ (
  .A(_057_),
  .B1(_097_),
  .B2(_172_),
  .ZN(_058_)
);

OAI21_X1 _291_ (
  .A(_056_),
  .B1(_058_),
  .B2(_100_),
  .ZN(_059_)
);

AOI21_X1 _292_ (
  .A(_118_),
  .B1(_055_),
  .B2(_059_),
  .ZN(_060_)
);

NAND3_X1 _293_ (
  .A1(_052_),
  .A2(_053_),
  .A3(_108_),
  .ZN(_061_)
);

NAND3_X1 _294_ (
  .A1(_061_),
  .A2(_111_),
  .A3(_027_),
  .ZN(_062_)
);

NOR2_X1 _295_ (
  .A1(_102_),
  .A2(_040_),
  .ZN(_063_)
);

OAI21_X1 _296_ (
  .A(_063_),
  .B1(_058_),
  .B2(_108_),
  .ZN(_064_)
);

NAND3_X1 _297_ (
  .A1(_062_),
  .A2(_064_),
  .A3(_120_),
  .ZN(_065_)
);

OAI21_X1 _298_ (
  .A(_051_),
  .B1(_060_),
  .B2(_065_),
  .ZN(_005_)
);

NAND2_X2 _299_ (
  .A1(_106_),
  .A2(_100_),
  .ZN(_066_)
);

NAND2_X1 _300_ (
  .A1(_099_),
  .A2(x[1]),
  .ZN(_067_)
);

NAND3_X1 _301_ (
  .A1(_066_),
  .A2(_103_),
  .A3(_067_),
  .ZN(_068_)
);

NAND2_X1 _302_ (
  .A1(_097_),
  .A2(_099_),
  .ZN(_069_)
);

OAI21_X1 _303_ (
  .A(_069_),
  .B1(_108_),
  .B2(x[1]),
  .ZN(_070_)
);

OAI21_X1 _304_ (
  .A(_068_),
  .B1(_070_),
  .B2(_103_),
  .ZN(_071_)
);

XNOR2_X1 _305_ (
  .A(_071_),
  .B(_116_),
  .ZN(_072_)
);

NAND2_X1 _306_ (
  .A1(_072_),
  .A2(_121_),
  .ZN(_073_)
);

NAND2_X1 _307_ (
  .A1(_123_),
  .A2(\coef[27] ),
  .ZN(_074_)
);

NAND2_X1 _308_ (
  .A1(_073_),
  .A2(_074_),
  .ZN(_006_)
);

NAND2_X1 _309_ (
  .A1(_047_),
  .A2(_040_),
  .ZN(_075_)
);

NAND2_X1 _310_ (
  .A1(_095_),
  .A2(_098_),
  .ZN(_076_)
);

OR2_X1 _311_ (
  .A1(_075_),
  .A2(_076_),
  .ZN(_077_)
);

NAND2_X1 _312_ (
  .A1(_075_),
  .A2(_076_),
  .ZN(_078_)
);

NAND3_X1 _313_ (
  .A1(_077_),
  .A2(_078_),
  .A3(_121_),
  .ZN(_079_)
);

INV_X1 _314_ (
  .A(\coef[28] ),
  .ZN(_080_)
);

OAI21_X1 _315_ (
  .A(_079_),
  .B1(_121_),
  .B2(_080_),
  .ZN(_007_)
);

NOR2_X1 _316_ (
  .A1(_121_),
  .A2(\coef[15] ),
  .ZN(_081_)
);

NAND2_X1 _317_ (
  .A1(_044_),
  .A2(_025_),
  .ZN(_082_)
);

NAND2_X1 _318_ (
  .A1(_082_),
  .A2(_027_),
  .ZN(_083_)
);

NAND2_X1 _319_ (
  .A1(_036_),
  .A2(_111_),
  .ZN(_084_)
);

NAND2_X1 _320_ (
  .A1(_084_),
  .A2(_031_),
  .ZN(_085_)
);

NAND2_X1 _321_ (
  .A1(_083_),
  .A2(_085_),
  .ZN(_086_)
);

AOI21_X1 _322_ (
  .A(_040_),
  .B1(_029_),
  .B2(_038_),
  .ZN(_087_)
);

NOR2_X1 _323_ (
  .A1(_086_),
  .A2(_087_),
  .ZN(_088_)
);

NAND2_X1 _324_ (
  .A1(_024_),
  .A2(_045_),
  .ZN(_089_)
);

AOI21_X1 _325_ (
  .A(_123_),
  .B1(_089_),
  .B2(_135_),
  .ZN(_090_)
);

AOI21_X2 _326_ (
  .A(_081_),
  .B1(_088_),
  .B2(_090_),
  .ZN(_008_)
);

NOR2_X1 _327_ (
  .A1(_121_),
  .A2(\coef[30] ),
  .ZN(_091_)
);

XNOR2_X1 _328_ (
  .A(_075_),
  .B(_093_),
  .ZN(_092_)
);

AOI21_X1 _329_ (
  .A(_091_),
  .B1(_092_),
  .B2(_121_),
  .ZN(_009_)
);

HA_X1 _330_ (
  .A(_160_),
  .B(_161_),
  .CO(_162_),
  .S(_163_)
);

HA_X1 _331_ (
  .A(_160_),
  .B(_161_),
  .CO(_164_),
  .S(_165_)
);

HA_X1 _332_ (
  .A(_160_),
  .B(x[1]),
  .CO(_166_),
  .S(_167_)
);

HA_X1 _333_ (
  .A(_160_),
  .B(x[1]),
  .CO(_168_),
  .S(_169_)
);

HA_X1 _334_ (
  .A(x[0]),
  .B(_161_),
  .CO(_170_),
  .S(_171_)
);

HA_X1 _335_ (
  .A(x[0]),
  .B(_161_),
  .CO(_172_),
  .S(_173_)
);

HA_X1 _336_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_174_),
  .S(_175_)
);

HA_X1 _337_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_176_),
  .S(_177_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_159_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_158_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_157_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_156_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_155_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_154_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_153_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_152_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_151_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_150_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$0c5a5bd6be4ed818deaac08b02afbddb6897ffee\dctu

module \$paramod$0f96740a02eb44c944b68d6b495a8cce162f1249\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _190_ (
  .A(x[1]),
  .ZN(_173_)
);

CLKBUF_X2 _191_ (
  .A(x[0]),
  .Z(_103_)
);

INV_X1 _192_ (
  .A(_103_),
  .ZN(_172_)
);

INV_X1 _193_ (
  .A(ena),
  .ZN(_104_)
);

BUF_X4 _194_ (
  .A(y[1]),
  .Z(_105_)
);

CLKBUF_X3 _195_ (
  .A(_105_),
  .Z(_106_)
);

BUF_X4 _196_ (
  .A(y[0]),
  .Z(_107_)
);

BUF_X4 _197_ (
  .A(_107_),
  .Z(_108_)
);

BUF_X4 _198_ (
  .A(x[2]),
  .Z(_109_)
);

INV_X8 _199_ (
  .A(_109_),
  .ZN(_110_)
);

BUF_X16 _200_ (
  .A(_110_),
  .Z(_111_)
);

INV_X1 _201_ (
  .A(_178_),
  .ZN(_112_)
);

NAND2_X2 _202_ (
  .A1(_111_),
  .A2(_112_),
  .ZN(_113_)
);

BUF_X8 _203_ (
  .A(_109_),
  .Z(_114_)
);

NAND2_X4 _204_ (
  .A1(_114_),
  .A2(_184_),
  .ZN(_115_)
);

AOI21_X2 _205_ (
  .A(_108_),
  .B1(_113_),
  .B2(_115_),
  .ZN(_116_)
);

INV_X4 _206_ (
  .A(_107_),
  .ZN(_117_)
);

NOR2_X1 _207_ (
  .A1(_117_),
  .A2(_103_),
  .ZN(_118_)
);

OAI21_X1 _208_ (
  .A(_106_),
  .B1(_116_),
  .B2(_118_),
  .ZN(_119_)
);

BUF_X1 _209_ (
  .A(y[2]),
  .Z(_120_)
);

INV_X1 _210_ (
  .A(_186_),
  .ZN(_121_)
);

NAND2_X4 _211_ (
  .A1(_111_),
  .A2(_121_),
  .ZN(_122_)
);

NAND2_X1 _212_ (
  .A1(_109_),
  .A2(_176_),
  .ZN(_123_)
);

NAND3_X1 _213_ (
  .A1(_122_),
  .A2(_108_),
  .A3(_123_),
  .ZN(_124_)
);

BUF_X8 _214_ (
  .A(_117_),
  .Z(_125_)
);

AOI21_X2 _215_ (
  .A(_105_),
  .B1(_125_),
  .B2(_114_),
  .ZN(_126_)
);

AOI21_X1 _216_ (
  .A(_120_),
  .B1(_124_),
  .B2(_126_),
  .ZN(_127_)
);

AOI21_X1 _217_ (
  .A(_104_),
  .B1(_119_),
  .B2(_127_),
  .ZN(_128_)
);

INV_X2 _218_ (
  .A(_105_),
  .ZN(_129_)
);

OR2_X1 _219_ (
  .A1(_180_),
  .A2(_109_),
  .ZN(_130_)
);

NAND2_X2 _220_ (
  .A1(_114_),
  .A2(_182_),
  .ZN(_131_)
);

NAND3_X1 _221_ (
  .A1(_130_),
  .A2(_108_),
  .A3(_131_),
  .ZN(_132_)
);

INV_X1 _222_ (
  .A(_132_),
  .ZN(_133_)
);

NOR2_X1 _223_ (
  .A1(_172_),
  .A2(_107_),
  .ZN(_134_)
);

OAI21_X1 _224_ (
  .A(_129_),
  .B1(_133_),
  .B2(_134_),
  .ZN(_135_)
);

INV_X1 _225_ (
  .A(_120_),
  .ZN(_136_)
);

INV_X1 _226_ (
  .A(_188_),
  .ZN(_137_)
);

NAND2_X4 _227_ (
  .A1(_111_),
  .A2(_137_),
  .ZN(_138_)
);

NAND2_X2 _228_ (
  .A1(_114_),
  .A2(_174_),
  .ZN(_139_)
);

NAND2_X1 _229_ (
  .A1(_138_),
  .A2(_139_),
  .ZN(_140_)
);

NAND2_X2 _230_ (
  .A1(_140_),
  .A2(_125_),
  .ZN(_141_)
);

NAND2_X4 _231_ (
  .A1(_111_),
  .A2(_107_),
  .ZN(_142_)
);

NAND2_X1 _232_ (
  .A1(_142_),
  .A2(_105_),
  .ZN(_143_)
);

INV_X1 _233_ (
  .A(_143_),
  .ZN(_144_)
);

AOI21_X1 _234_ (
  .A(_136_),
  .B1(_141_),
  .B2(_144_),
  .ZN(_145_)
);

NAND2_X1 _235_ (
  .A1(_135_),
  .A2(_145_),
  .ZN(_146_)
);

NAND2_X1 _236_ (
  .A1(_128_),
  .A2(_146_),
  .ZN(_147_)
);

NAND2_X1 _237_ (
  .A1(_104_),
  .A2(\coef[21] ),
  .ZN(_148_)
);

NAND2_X1 _238_ (
  .A1(_147_),
  .A2(_148_),
  .ZN(_000_)
);

NAND2_X2 _239_ (
  .A1(_117_),
  .A2(_114_),
  .ZN(_149_)
);

NAND2_X1 _240_ (
  .A1(_117_),
  .A2(_172_),
  .ZN(_150_)
);

MUX2_X1 _241_ (
  .A(_149_),
  .B(_150_),
  .S(_105_),
  .Z(_151_)
);

NAND3_X2 _242_ (
  .A1(_138_),
  .A2(_107_),
  .A3(_139_),
  .ZN(_152_)
);

NAND3_X1 _243_ (
  .A1(_151_),
  .A2(_136_),
  .A3(_152_),
  .ZN(_153_)
);

BUF_X2 _244_ (
  .A(ena),
  .Z(_154_)
);

NAND2_X1 _245_ (
  .A1(_108_),
  .A2(_103_),
  .ZN(_155_)
);

INV_X1 _246_ (
  .A(_155_),
  .ZN(_156_)
);

OAI21_X1 _247_ (
  .A(_143_),
  .B1(_106_),
  .B2(_156_),
  .ZN(_157_)
);

NAND2_X4 _248_ (
  .A1(_122_),
  .A2(_123_),
  .ZN(_158_)
);

NAND2_X4 _249_ (
  .A1(_158_),
  .A2(_125_),
  .ZN(_159_)
);

BUF_X2 _250_ (
  .A(_120_),
  .Z(_160_)
);

NAND3_X1 _251_ (
  .A1(_157_),
  .A2(_159_),
  .A3(_160_),
  .ZN(_161_)
);

NAND3_X1 _252_ (
  .A1(_153_),
  .A2(_154_),
  .A3(_161_),
  .ZN(_162_)
);

NAND2_X1 _253_ (
  .A1(_104_),
  .A2(\coef[23] ),
  .ZN(_009_)
);

NAND2_X1 _254_ (
  .A1(_162_),
  .A2(_009_),
  .ZN(_001_)
);

INV_X1 _255_ (
  .A(_182_),
  .ZN(_010_)
);

NAND2_X4 _256_ (
  .A1(_111_),
  .A2(_010_),
  .ZN(_011_)
);

NAND2_X1 _257_ (
  .A1(_109_),
  .A2(_180_),
  .ZN(_012_)
);

NAND2_X2 _258_ (
  .A1(_011_),
  .A2(_012_),
  .ZN(_013_)
);

NAND2_X2 _259_ (
  .A1(_013_),
  .A2(_108_),
  .ZN(_014_)
);

NAND2_X1 _260_ (
  .A1(_159_),
  .A2(_014_),
  .ZN(_015_)
);

NAND2_X1 _261_ (
  .A1(_015_),
  .A2(_106_),
  .ZN(_016_)
);

INV_X1 _262_ (
  .A(_134_),
  .ZN(_017_)
);

NAND2_X1 _263_ (
  .A1(_108_),
  .A2(x[1]),
  .ZN(_018_)
);

NAND3_X1 _264_ (
  .A1(_017_),
  .A2(_018_),
  .A3(_129_),
  .ZN(_019_)
);

NAND3_X1 _265_ (
  .A1(_016_),
  .A2(_160_),
  .A3(_019_),
  .ZN(_020_)
);

NOR2_X1 _266_ (
  .A1(_107_),
  .A2(x[1]),
  .ZN(_021_)
);

NOR3_X1 _267_ (
  .A1(_118_),
  .A2(_021_),
  .A3(_129_),
  .ZN(_022_)
);

NOR2_X1 _268_ (
  .A1(_022_),
  .A2(_160_),
  .ZN(_023_)
);

NAND2_X1 _269_ (
  .A1(_110_),
  .A2(_184_),
  .ZN(_024_)
);

NAND2_X1 _270_ (
  .A1(_112_),
  .A2(_109_),
  .ZN(_025_)
);

NAND2_X1 _271_ (
  .A1(_024_),
  .A2(_025_),
  .ZN(_026_)
);

NAND2_X2 _272_ (
  .A1(_026_),
  .A2(_125_),
  .ZN(_027_)
);

NAND2_X1 _273_ (
  .A1(_027_),
  .A2(_152_),
  .ZN(_028_)
);

NAND2_X1 _274_ (
  .A1(_028_),
  .A2(_129_),
  .ZN(_029_)
);

NAND2_X1 _275_ (
  .A1(_023_),
  .A2(_029_),
  .ZN(_030_)
);

NAND3_X1 _276_ (
  .A1(_020_),
  .A2(_154_),
  .A3(_030_),
  .ZN(_031_)
);

NAND2_X1 _277_ (
  .A1(_104_),
  .A2(\coef[24] ),
  .ZN(_032_)
);

NAND2_X1 _278_ (
  .A1(_031_),
  .A2(_032_),
  .ZN(_002_)
);

NAND2_X1 _279_ (
  .A1(_111_),
  .A2(_174_),
  .ZN(_033_)
);

NAND2_X1 _280_ (
  .A1(_137_),
  .A2(_114_),
  .ZN(_034_)
);

NAND3_X1 _281_ (
  .A1(_033_),
  .A2(_034_),
  .A3(_108_),
  .ZN(_035_)
);

NAND2_X1 _282_ (
  .A1(_027_),
  .A2(_035_),
  .ZN(_036_)
);

NAND2_X1 _283_ (
  .A1(_036_),
  .A2(_129_),
  .ZN(_037_)
);

NAND2_X1 _284_ (
  .A1(_111_),
  .A2(_180_),
  .ZN(_038_)
);

NAND2_X1 _285_ (
  .A1(_010_),
  .A2(_114_),
  .ZN(_039_)
);

NAND3_X1 _286_ (
  .A1(_038_),
  .A2(_039_),
  .A3(_125_),
  .ZN(_040_)
);

NAND3_X1 _287_ (
  .A1(_040_),
  .A2(_124_),
  .A3(_106_),
  .ZN(_041_)
);

NAND3_X1 _288_ (
  .A1(_037_),
  .A2(_041_),
  .A3(_160_),
  .ZN(_042_)
);

INV_X1 _289_ (
  .A(_176_),
  .ZN(_043_)
);

NAND2_X2 _290_ (
  .A1(_111_),
  .A2(_043_),
  .ZN(_044_)
);

NAND2_X1 _291_ (
  .A1(_114_),
  .A2(_186_),
  .ZN(_045_)
);

NAND3_X1 _292_ (
  .A1(_044_),
  .A2(_125_),
  .A3(_045_),
  .ZN(_046_)
);

NAND2_X1 _293_ (
  .A1(_014_),
  .A2(_046_),
  .ZN(_047_)
);

NAND2_X1 _294_ (
  .A1(_047_),
  .A2(_106_),
  .ZN(_048_)
);

NAND3_X1 _295_ (
  .A1(_113_),
  .A2(_108_),
  .A3(_115_),
  .ZN(_049_)
);

NAND3_X1 _296_ (
  .A1(_141_),
  .A2(_049_),
  .A3(_129_),
  .ZN(_050_)
);

NAND3_X1 _297_ (
  .A1(_048_),
  .A2(_050_),
  .A3(_136_),
  .ZN(_051_)
);

NAND3_X1 _298_ (
  .A1(_042_),
  .A2(_051_),
  .A3(_154_),
  .ZN(_052_)
);

NAND2_X1 _299_ (
  .A1(_104_),
  .A2(\coef[10] ),
  .ZN(_053_)
);

NAND2_X1 _300_ (
  .A1(_052_),
  .A2(_053_),
  .ZN(_003_)
);

NAND2_X1 _301_ (
  .A1(_149_),
  .A2(_105_),
  .ZN(_054_)
);

INV_X1 _302_ (
  .A(_054_),
  .ZN(_055_)
);

AOI21_X1 _303_ (
  .A(_120_),
  .B1(_055_),
  .B2(_142_),
  .ZN(_056_)
);

NAND2_X1 _304_ (
  .A1(_132_),
  .A2(_159_),
  .ZN(_057_)
);

INV_X1 _305_ (
  .A(_057_),
  .ZN(_058_)
);

OAI21_X2 _306_ (
  .A(_056_),
  .B1(_058_),
  .B2(_106_),
  .ZN(_059_)
);

INV_X1 _307_ (
  .A(_152_),
  .ZN(_060_)
);

OAI21_X1 _308_ (
  .A(_106_),
  .B1(_060_),
  .B2(_116_),
  .ZN(_061_)
);

AOI21_X1 _309_ (
  .A(_136_),
  .B1(_126_),
  .B2(_142_),
  .ZN(_062_)
);

NAND2_X1 _310_ (
  .A1(_061_),
  .A2(_062_),
  .ZN(_063_)
);

NAND3_X1 _311_ (
  .A1(_059_),
  .A2(_063_),
  .A3(_154_),
  .ZN(_064_)
);

NAND2_X1 _312_ (
  .A1(_104_),
  .A2(\coef[26] ),
  .ZN(_065_)
);

NAND2_X1 _313_ (
  .A1(_064_),
  .A2(_065_),
  .ZN(_004_)
);

NOR2_X1 _314_ (
  .A1(_154_),
  .A2(\coef[13] ),
  .ZN(_066_)
);

NOR2_X1 _315_ (
  .A1(_021_),
  .A2(_105_),
  .ZN(_067_)
);

AOI21_X1 _316_ (
  .A(_160_),
  .B1(_014_),
  .B2(_067_),
  .ZN(_068_)
);

NAND3_X1 _317_ (
  .A1(_033_),
  .A2(_034_),
  .A3(_125_),
  .ZN(_069_)
);

INV_X1 _318_ (
  .A(_175_),
  .ZN(_070_)
);

NAND2_X4 _319_ (
  .A1(_111_),
  .A2(_070_),
  .ZN(_071_)
);

NAND2_X4 _320_ (
  .A1(_114_),
  .A2(_175_),
  .ZN(_072_)
);

NAND3_X2 _321_ (
  .A1(_071_),
  .A2(_108_),
  .A3(_072_),
  .ZN(_073_)
);

NAND3_X1 _322_ (
  .A1(_069_),
  .A2(_073_),
  .A3(_106_),
  .ZN(_074_)
);

AOI21_X1 _323_ (
  .A(_104_),
  .B1(_068_),
  .B2(_074_),
  .ZN(_075_)
);

NAND2_X2 _324_ (
  .A1(_071_),
  .A2(_072_),
  .ZN(_076_)
);

NAND2_X2 _325_ (
  .A1(_076_),
  .A2(_125_),
  .ZN(_077_)
);

NAND3_X1 _326_ (
  .A1(_044_),
  .A2(_108_),
  .A3(_045_),
  .ZN(_078_)
);

NAND3_X1 _327_ (
  .A1(_077_),
  .A2(_078_),
  .A3(_129_),
  .ZN(_079_)
);

NAND3_X1 _328_ (
  .A1(_027_),
  .A2(_106_),
  .A3(_018_),
  .ZN(_080_)
);

NAND3_X1 _329_ (
  .A1(_079_),
  .A2(_080_),
  .A3(_160_),
  .ZN(_081_)
);

AOI21_X1 _330_ (
  .A(_066_),
  .B1(_075_),
  .B2(_081_),
  .ZN(_005_)
);

NAND3_X1 _331_ (
  .A1(_077_),
  .A2(_129_),
  .A3(_142_),
  .ZN(_082_)
);

NAND2_X1 _332_ (
  .A1(_023_),
  .A2(_082_),
  .ZN(_083_)
);

NAND2_X1 _333_ (
  .A1(_073_),
  .A2(_055_),
  .ZN(_084_)
);

NAND3_X1 _334_ (
  .A1(_084_),
  .A2(_160_),
  .A3(_019_),
  .ZN(_085_)
);

NAND3_X1 _335_ (
  .A1(_083_),
  .A2(_154_),
  .A3(_085_),
  .ZN(_086_)
);

INV_X1 _336_ (
  .A(\coef[28] ),
  .ZN(_087_)
);

OAI21_X1 _337_ (
  .A(_086_),
  .B1(_154_),
  .B2(_087_),
  .ZN(_006_)
);

NAND2_X1 _338_ (
  .A1(_104_),
  .A2(\coef[29] ),
  .ZN(_088_)
);

NAND3_X1 _339_ (
  .A1(_071_),
  .A2(_125_),
  .A3(_072_),
  .ZN(_089_)
);

NAND3_X1 _340_ (
  .A1(_049_),
  .A2(_089_),
  .A3(_105_),
  .ZN(_090_)
);

NAND3_X1 _341_ (
  .A1(_010_),
  .A2(_111_),
  .A3(_107_),
  .ZN(_091_)
);

NAND3_X1 _342_ (
  .A1(_114_),
  .A2(_107_),
  .A3(_180_),
  .ZN(_092_)
);

NAND3_X1 _343_ (
  .A1(_091_),
  .A2(_092_),
  .A3(_150_),
  .ZN(_093_)
);

NAND2_X1 _344_ (
  .A1(_093_),
  .A2(_129_),
  .ZN(_094_)
);

NAND3_X1 _345_ (
  .A1(_090_),
  .A2(_094_),
  .A3(_160_),
  .ZN(_095_)
);

NAND2_X1 _346_ (
  .A1(_095_),
  .A2(_154_),
  .ZN(_096_)
);

NAND3_X1 _347_ (
  .A1(_130_),
  .A2(_125_),
  .A3(_131_),
  .ZN(_097_)
);

NAND3_X1 _348_ (
  .A1(_097_),
  .A2(_073_),
  .A3(_129_),
  .ZN(_098_)
);

NAND3_X1 _349_ (
  .A1(_027_),
  .A2(_106_),
  .A3(_155_),
  .ZN(_099_)
);

AOI21_X1 _350_ (
  .A(_160_),
  .B1(_098_),
  .B2(_099_),
  .ZN(_100_)
);

OAI21_X1 _351_ (
  .A(_088_),
  .B1(_096_),
  .B2(_100_),
  .ZN(_007_)
);

NOR2_X1 _352_ (
  .A1(_154_),
  .A2(\coef[30] ),
  .ZN(_101_)
);

XNOR2_X1 _353_ (
  .A(_160_),
  .B(_103_),
  .ZN(_102_)
);

AOI21_X1 _354_ (
  .A(_101_),
  .B1(_102_),
  .B2(_154_),
  .ZN(_008_)
);

HA_X1 _355_ (
  .A(_172_),
  .B(_173_),
  .CO(_174_),
  .S(_175_)
);

HA_X1 _356_ (
  .A(_172_),
  .B(_173_),
  .CO(_176_),
  .S(_177_)
);

HA_X1 _357_ (
  .A(_172_),
  .B(x[1]),
  .CO(_178_),
  .S(_179_)
);

HA_X1 _358_ (
  .A(_172_),
  .B(x[1]),
  .CO(_180_),
  .S(_181_)
);

HA_X1 _359_ (
  .A(x[0]),
  .B(_173_),
  .CO(_182_),
  .S(_183_)
);

HA_X1 _360_ (
  .A(x[0]),
  .B(_173_),
  .CO(_184_),
  .S(_185_)
);

HA_X1 _361_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_186_),
  .S(_187_)
);

HA_X1 _362_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_188_),
  .S(_189_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_171_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_170_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_169_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_168_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_167_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_166_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_165_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_164_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_163_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$0f96740a02eb44c944b68d6b495a8cce162f1249\dctu

module \$paramod$88a8287894fa5d106cca0ce24429339f4a2785a9\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X2 _054_ (
  .A(x[2]),
  .ZN(_004_)
);

INV_X1 _055_ (
  .A(x[0]),
  .ZN(_005_)
);

NAND2_X2 _056_ (
  .A1(_004_),
  .A2(_005_),
  .ZN(_006_)
);

NAND2_X1 _057_ (
  .A1(x[2]),
  .A2(x[0]),
  .ZN(_007_)
);

NAND2_X2 _058_ (
  .A1(_006_),
  .A2(_007_),
  .ZN(_008_)
);

NAND2_X2 _059_ (
  .A1(_008_),
  .A2(y[0]),
  .ZN(_009_)
);

INV_X1 _060_ (
  .A(x[1]),
  .ZN(_010_)
);

NAND2_X1 _061_ (
  .A1(_004_),
  .A2(_010_),
  .ZN(_011_)
);

INV_X1 _062_ (
  .A(y[0]),
  .ZN(_012_)
);

NAND2_X1 _063_ (
  .A1(x[2]),
  .A2(x[1]),
  .ZN(_013_)
);

NAND3_X1 _064_ (
  .A1(_011_),
  .A2(_012_),
  .A3(_013_),
  .ZN(_014_)
);

NAND2_X1 _065_ (
  .A1(_009_),
  .A2(_014_),
  .ZN(_015_)
);

CLKBUF_X2 _066_ (
  .A(y[1]),
  .Z(_016_)
);

NAND2_X1 _067_ (
  .A1(_015_),
  .A2(_016_),
  .ZN(_017_)
);

NAND2_X1 _068_ (
  .A1(_011_),
  .A2(_013_),
  .ZN(_018_)
);

NAND2_X2 _069_ (
  .A1(_018_),
  .A2(y[0]),
  .ZN(_019_)
);

NAND3_X1 _070_ (
  .A1(_006_),
  .A2(_012_),
  .A3(_007_),
  .ZN(_020_)
);

NAND2_X1 _071_ (
  .A1(_019_),
  .A2(_020_),
  .ZN(_021_)
);

INV_X1 _072_ (
  .A(_016_),
  .ZN(_022_)
);

NAND2_X1 _073_ (
  .A1(_021_),
  .A2(_022_),
  .ZN(_023_)
);

BUF_X1 _074_ (
  .A(y[2]),
  .Z(_024_)
);

INV_X1 _075_ (
  .A(_024_),
  .ZN(_025_)
);

NAND3_X1 _076_ (
  .A1(_017_),
  .A2(_023_),
  .A3(_025_),
  .ZN(_026_)
);

NAND3_X1 _077_ (
  .A1(_019_),
  .A2(_020_),
  .A3(_022_),
  .ZN(_027_)
);

NAND3_X1 _078_ (
  .A1(_009_),
  .A2(_014_),
  .A3(_016_),
  .ZN(_028_)
);

NAND3_X1 _079_ (
  .A1(_027_),
  .A2(_028_),
  .A3(_024_),
  .ZN(_029_)
);

BUF_X2 _080_ (
  .A(ena),
  .Z(_030_)
);

NAND3_X1 _081_ (
  .A1(_026_),
  .A2(_029_),
  .A3(_030_),
  .ZN(_031_)
);

INV_X1 _082_ (
  .A(_030_),
  .ZN(_032_)
);

NAND2_X1 _083_ (
  .A1(_032_),
  .A2(\coef[13] ),
  .ZN(_033_)
);

NAND2_X1 _084_ (
  .A1(_031_),
  .A2(_033_),
  .ZN(_000_)
);

NAND3_X1 _085_ (
  .A1(_017_),
  .A2(_023_),
  .A3(_024_),
  .ZN(_034_)
);

NAND3_X1 _086_ (
  .A1(_027_),
  .A2(_028_),
  .A3(_025_),
  .ZN(_035_)
);

NAND3_X1 _087_ (
  .A1(_034_),
  .A2(_035_),
  .A3(_030_),
  .ZN(_036_)
);

NAND2_X1 _088_ (
  .A1(_032_),
  .A2(\coef[10] ),
  .ZN(_037_)
);

NAND2_X1 _089_ (
  .A1(_036_),
  .A2(_037_),
  .ZN(_001_)
);

NAND2_X1 _090_ (
  .A1(_008_),
  .A2(_012_),
  .ZN(_038_)
);

NAND3_X1 _091_ (
  .A1(_038_),
  .A2(_019_),
  .A3(_016_),
  .ZN(_039_)
);

NAND3_X1 _092_ (
  .A1(_006_),
  .A2(y[0]),
  .A3(_007_),
  .ZN(_040_)
);

NAND3_X1 _093_ (
  .A1(_040_),
  .A2(_014_),
  .A3(_022_),
  .ZN(_041_)
);

NAND2_X1 _094_ (
  .A1(_039_),
  .A2(_041_),
  .ZN(_042_)
);

NAND2_X1 _095_ (
  .A1(_042_),
  .A2(_025_),
  .ZN(_043_)
);

NAND3_X1 _096_ (
  .A1(_039_),
  .A2(_041_),
  .A3(_024_),
  .ZN(_044_)
);

NAND3_X1 _097_ (
  .A1(_043_),
  .A2(_044_),
  .A3(_030_),
  .ZN(_045_)
);

NAND2_X1 _098_ (
  .A1(_032_),
  .A2(\coef[29] ),
  .ZN(_046_)
);

NAND2_X1 _099_ (
  .A1(_045_),
  .A2(_046_),
  .ZN(_002_)
);

NOR2_X1 _100_ (
  .A1(_030_),
  .A2(\coef[30] ),
  .ZN(_047_)
);

XNOR2_X1 _101_ (
  .A(_016_),
  .B(_024_),
  .ZN(_048_)
);

XNOR2_X1 _102_ (
  .A(_048_),
  .B(_008_),
  .ZN(_049_)
);

AOI21_X1 _103_ (
  .A(_047_),
  .B1(_049_),
  .B2(_030_),
  .ZN(_003_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_053_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_052_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_051_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_050_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[10] , \coef[13] , \coef[10] , \coef[10] , \coef[13] , \coef[10] , \coef[13] , \coef[10] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$88a8287894fa5d106cca0ce24429339f4a2785a9\dctu

module \$paramod$8cd9bf70556f3aa976ca66d64ee3b9c1b3a94e21\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _0_;
wire _1_;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_85002  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({_1_, _1_, _0_, _1_, _1_, _1_, _1_, _1_, _1_, _1_, _1_}),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$8cd9bf70556f3aa976ca66d64ee3b9c1b3a94e21\dctu

module \$paramod$8f6708f3156f3d6d195809cddd67c9b8c08cd488\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X2 _066_ (
  .A(x[1]),
  .ZN(_008_)
);

NAND2_X2 _067_ (
  .A1(_008_),
  .A2(x[0]),
  .ZN(_009_)
);

INV_X2 _068_ (
  .A(x[0]),
  .ZN(_010_)
);

NAND2_X2 _069_ (
  .A1(_010_),
  .A2(x[1]),
  .ZN(_011_)
);

NAND3_X4 _070_ (
  .A1(_009_),
  .A2(_011_),
  .A3(y[0]),
  .ZN(_012_)
);

NAND2_X2 _071_ (
  .A1(_008_),
  .A2(_010_),
  .ZN(_013_)
);

INV_X1 _072_ (
  .A(y[0]),
  .ZN(_014_)
);

NAND2_X1 _073_ (
  .A1(x[1]),
  .A2(x[0]),
  .ZN(_015_)
);

NAND3_X4 _074_ (
  .A1(_013_),
  .A2(_014_),
  .A3(_015_),
  .ZN(_016_)
);

NAND2_X4 _075_ (
  .A1(_012_),
  .A2(_016_),
  .ZN(_017_)
);

NAND2_X2 _076_ (
  .A1(_017_),
  .A2(y[1]),
  .ZN(_018_)
);

NAND2_X2 _077_ (
  .A1(_009_),
  .A2(_011_),
  .ZN(_019_)
);

INV_X1 _078_ (
  .A(y[1]),
  .ZN(_020_)
);

NAND2_X1 _079_ (
  .A1(_019_),
  .A2(_020_),
  .ZN(_021_)
);

BUF_X4 _080_ (
  .A(ena),
  .Z(_022_)
);

INV_X2 _081_ (
  .A(_022_),
  .ZN(_023_)
);

BUF_X1 _082_ (
  .A(y[2]),
  .Z(_024_)
);

NOR2_X1 _083_ (
  .A1(_023_),
  .A2(_024_),
  .ZN(_025_)
);

NAND3_X1 _084_ (
  .A1(_018_),
  .A2(_021_),
  .A3(_025_),
  .ZN(_026_)
);

NAND3_X1 _085_ (
  .A1(_009_),
  .A2(_011_),
  .A3(_014_),
  .ZN(_027_)
);

NAND3_X1 _086_ (
  .A1(_013_),
  .A2(y[0]),
  .A3(_015_),
  .ZN(_028_)
);

NAND3_X1 _087_ (
  .A1(_027_),
  .A2(_028_),
  .A3(_020_),
  .ZN(_029_)
);

NOR2_X2 _088_ (
  .A1(_019_),
  .A2(_020_),
  .ZN(_030_)
);

NOR2_X2 _089_ (
  .A1(_030_),
  .A2(_023_),
  .ZN(_031_)
);

NAND3_X1 _090_ (
  .A1(_029_),
  .A2(_024_),
  .A3(_031_),
  .ZN(_032_)
);

NAND2_X1 _091_ (
  .A1(_023_),
  .A2(\coef[21] ),
  .ZN(_033_)
);

NAND3_X1 _092_ (
  .A1(_026_),
  .A2(_032_),
  .A3(_033_),
  .ZN(_000_)
);

NAND3_X2 _093_ (
  .A1(_012_),
  .A2(_016_),
  .A3(_020_),
  .ZN(_034_)
);

INV_X1 _094_ (
  .A(_024_),
  .ZN(_035_)
);

NAND3_X1 _095_ (
  .A1(_018_),
  .A2(_034_),
  .A3(_035_),
  .ZN(_036_)
);

NAND3_X2 _096_ (
  .A1(_012_),
  .A2(_016_),
  .A3(y[1]),
  .ZN(_037_)
);

NAND3_X1 _097_ (
  .A1(_037_),
  .A2(_029_),
  .A3(_024_),
  .ZN(_038_)
);

NAND3_X1 _098_ (
  .A1(_036_),
  .A2(_038_),
  .A3(_022_),
  .ZN(_039_)
);

NAND2_X1 _099_ (
  .A1(_023_),
  .A2(\coef[22] ),
  .ZN(_040_)
);

NAND2_X1 _100_ (
  .A1(_039_),
  .A2(_040_),
  .ZN(_001_)
);

MUX2_X1 _101_ (
  .A(\coef[23] ),
  .B(_017_),
  .S(_022_),
  .Z(_002_)
);

NAND3_X1 _102_ (
  .A1(_037_),
  .A2(_029_),
  .A3(_035_),
  .ZN(_041_)
);

NAND3_X1 _103_ (
  .A1(_018_),
  .A2(_034_),
  .A3(_024_),
  .ZN(_042_)
);

NAND3_X1 _104_ (
  .A1(_041_),
  .A2(_042_),
  .A3(_022_),
  .ZN(_043_)
);

NAND2_X1 _105_ (
  .A1(_023_),
  .A2(\coef[14] ),
  .ZN(_044_)
);

NAND2_X1 _106_ (
  .A1(_043_),
  .A2(_044_),
  .ZN(_003_)
);

NAND2_X1 _107_ (
  .A1(_037_),
  .A2(_021_),
  .ZN(_045_)
);

NAND3_X1 _108_ (
  .A1(_045_),
  .A2(_024_),
  .A3(_022_),
  .ZN(_046_)
);

INV_X2 _109_ (
  .A(_034_),
  .ZN(_047_)
);

OAI21_X1 _110_ (
  .A(_025_),
  .B1(_047_),
  .B2(_030_),
  .ZN(_048_)
);

NAND2_X1 _111_ (
  .A1(_023_),
  .A2(\coef[13] ),
  .ZN(_049_)
);

NAND3_X1 _112_ (
  .A1(_046_),
  .A2(_048_),
  .A3(_049_),
  .ZN(_004_)
);

NAND3_X1 _113_ (
  .A1(_037_),
  .A2(_021_),
  .A3(_025_),
  .ZN(_050_)
);

OAI21_X1 _114_ (
  .A(_050_),
  .B1(_022_),
  .B2(\coef[28] ),
  .ZN(_051_)
);

NAND2_X1 _115_ (
  .A1(_024_),
  .A2(_022_),
  .ZN(_052_)
);

NOR3_X2 _116_ (
  .A1(_047_),
  .A2(_030_),
  .A3(_052_),
  .ZN(_053_)
);

NOR2_X2 _117_ (
  .A1(_051_),
  .A2(_053_),
  .ZN(_005_)
);

NAND2_X1 _118_ (
  .A1(_031_),
  .A2(_021_),
  .ZN(_054_)
);

INV_X1 _119_ (
  .A(\coef[15] ),
  .ZN(_055_)
);

OAI21_X1 _120_ (
  .A(_054_),
  .B1(_022_),
  .B2(_055_),
  .ZN(_006_)
);

INV_X1 _121_ (
  .A(_019_),
  .ZN(_056_)
);

OAI22_X1 _122_ (
  .A1(_056_),
  .A2(_052_),
  .B1(\coef[12] ),
  .B2(_022_),
  .ZN(_057_)
);

AOI21_X1 _123_ (
  .A(_057_),
  .B1(_025_),
  .B2(_056_),
  .ZN(_007_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_065_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_064_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_063_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_062_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_061_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_060_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_059_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_058_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$8f6708f3156f3d6d195809cddd67c9b8c08cd488\dctu

module \$paramod$94a1b10314722615b96d6c8f661cbb82ecebf320\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _175_ (
  .A(x[0]),
  .ZN(_157_)
);

INV_X1 _176_ (
  .A(x[1]),
  .ZN(_158_)
);

BUF_X8 _177_ (
  .A(x[2]),
  .Z(_090_)
);

INV_X8 _178_ (
  .A(_090_),
  .ZN(_091_)
);

INV_X1 _179_ (
  .A(_160_),
  .ZN(_092_)
);

NAND2_X4 _180_ (
  .A1(_091_),
  .A2(_092_),
  .ZN(_093_)
);

NAND2_X4 _181_ (
  .A1(_090_),
  .A2(_160_),
  .ZN(_094_)
);

NAND2_X4 _182_ (
  .A1(_093_),
  .A2(_094_),
  .ZN(_095_)
);

BUF_X4 _183_ (
  .A(y[0]),
  .Z(_096_)
);

BUF_X8 _184_ (
  .A(_096_),
  .Z(_097_)
);

NAND2_X4 _185_ (
  .A1(_095_),
  .A2(_097_),
  .ZN(_098_)
);

NOR2_X2 _186_ (
  .A1(_157_),
  .A2(_096_),
  .ZN(_099_)
);

BUF_X4 _187_ (
  .A(y[1]),
  .Z(_100_)
);

NOR2_X2 _188_ (
  .A1(_099_),
  .A2(_100_),
  .ZN(_101_)
);

NAND2_X2 _189_ (
  .A1(_098_),
  .A2(_101_),
  .ZN(_102_)
);

INV_X8 _190_ (
  .A(_096_),
  .ZN(_103_)
);

NAND3_X4 _191_ (
  .A1(_093_),
  .A2(_103_),
  .A3(_094_),
  .ZN(_104_)
);

OAI21_X2 _192_ (
  .A(_100_),
  .B1(_103_),
  .B2(x[0]),
  .ZN(_105_)
);

INV_X1 _193_ (
  .A(_105_),
  .ZN(_106_)
);

NAND2_X2 _194_ (
  .A1(_104_),
  .A2(_106_),
  .ZN(_107_)
);

NAND2_X1 _195_ (
  .A1(_102_),
  .A2(_107_),
  .ZN(_108_)
);

BUF_X4 _196_ (
  .A(y[2]),
  .Z(_109_)
);

INV_X4 _197_ (
  .A(_109_),
  .ZN(_110_)
);

NAND2_X1 _198_ (
  .A1(_108_),
  .A2(_110_),
  .ZN(_111_)
);

NAND3_X1 _199_ (
  .A1(_102_),
  .A2(_107_),
  .A3(_109_),
  .ZN(_112_)
);

BUF_X2 _200_ (
  .A(ena),
  .Z(_113_)
);

BUF_X4 _201_ (
  .A(_113_),
  .Z(_114_)
);

NAND3_X1 _202_ (
  .A1(_111_),
  .A2(_112_),
  .A3(_114_),
  .ZN(_115_)
);

INV_X1 _203_ (
  .A(_113_),
  .ZN(_116_)
);

NAND2_X1 _204_ (
  .A1(_116_),
  .A2(\coef[21] ),
  .ZN(_117_)
);

NAND2_X1 _205_ (
  .A1(_115_),
  .A2(_117_),
  .ZN(_000_)
);

NOR2_X1 _206_ (
  .A1(_113_),
  .A2(\coef[22] ),
  .ZN(_118_)
);

NOR2_X2 _207_ (
  .A1(_110_),
  .A2(_100_),
  .ZN(_119_)
);

INV_X4 _208_ (
  .A(_100_),
  .ZN(_120_)
);

NOR2_X4 _209_ (
  .A1(_120_),
  .A2(_109_),
  .ZN(_121_)
);

NOR2_X2 _210_ (
  .A1(_119_),
  .A2(_121_),
  .ZN(_122_)
);

BUF_X16 _211_ (
  .A(_090_),
  .Z(_123_)
);

XNOR2_X1 _212_ (
  .A(_122_),
  .B(_123_),
  .ZN(_124_)
);

AOI21_X1 _213_ (
  .A(_118_),
  .B1(_124_),
  .B2(_114_),
  .ZN(_001_)
);

NAND2_X1 _214_ (
  .A1(_116_),
  .A2(\coef[23] ),
  .ZN(_125_)
);

INV_X1 _215_ (
  .A(_159_),
  .ZN(_126_)
);

NAND2_X1 _216_ (
  .A1(_091_),
  .A2(_126_),
  .ZN(_127_)
);

NAND2_X4 _217_ (
  .A1(_123_),
  .A2(_173_),
  .ZN(_128_)
);

NAND2_X1 _218_ (
  .A1(_127_),
  .A2(_128_),
  .ZN(_129_)
);

NAND2_X1 _219_ (
  .A1(_129_),
  .A2(_103_),
  .ZN(_130_)
);

NAND2_X1 _220_ (
  .A1(_100_),
  .A2(_109_),
  .ZN(_131_)
);

INV_X1 _221_ (
  .A(_131_),
  .ZN(_132_)
);

NAND3_X1 _222_ (
  .A1(_098_),
  .A2(_130_),
  .A3(_132_),
  .ZN(_133_)
);

NAND3_X1 _223_ (
  .A1(_127_),
  .A2(_097_),
  .A3(_128_),
  .ZN(_134_)
);

NAND2_X1 _224_ (
  .A1(_104_),
  .A2(_134_),
  .ZN(_135_)
);

NOR2_X1 _225_ (
  .A1(_100_),
  .A2(_109_),
  .ZN(_136_)
);

NAND2_X1 _226_ (
  .A1(_135_),
  .A2(_136_),
  .ZN(_137_)
);

INV_X1 _227_ (
  .A(_161_),
  .ZN(_138_)
);

NAND2_X1 _228_ (
  .A1(_091_),
  .A2(_138_),
  .ZN(_139_)
);

NAND2_X1 _229_ (
  .A1(_123_),
  .A2(_171_),
  .ZN(_140_)
);

NAND3_X1 _230_ (
  .A1(_139_),
  .A2(_103_),
  .A3(_140_),
  .ZN(_141_)
);

NAND3_X1 _231_ (
  .A1(_093_),
  .A2(_097_),
  .A3(_094_),
  .ZN(_142_)
);

NAND3_X1 _232_ (
  .A1(_141_),
  .A2(_142_),
  .A3(_121_),
  .ZN(_143_)
);

NAND3_X1 _233_ (
  .A1(_133_),
  .A2(_137_),
  .A3(_143_),
  .ZN(_144_)
);

NAND3_X1 _234_ (
  .A1(_139_),
  .A2(_097_),
  .A3(_140_),
  .ZN(_145_)
);

NAND3_X1 _235_ (
  .A1(_145_),
  .A2(_104_),
  .A3(_119_),
  .ZN(_146_)
);

NAND2_X1 _236_ (
  .A1(_146_),
  .A2(_114_),
  .ZN(_010_)
);

OAI21_X2 _237_ (
  .A(_125_),
  .B1(_144_),
  .B2(_010_),
  .ZN(_002_)
);

NAND2_X1 _238_ (
  .A1(_116_),
  .A2(\coef[24] ),
  .ZN(_011_)
);

NAND2_X1 _239_ (
  .A1(_126_),
  .A2(_123_),
  .ZN(_012_)
);

NAND2_X1 _240_ (
  .A1(_091_),
  .A2(_173_),
  .ZN(_013_)
);

NAND3_X1 _241_ (
  .A1(_122_),
  .A2(_012_),
  .A3(_013_),
  .ZN(_014_)
);

NAND2_X1 _242_ (
  .A1(_014_),
  .A2(_114_),
  .ZN(_015_)
);

NAND2_X1 _243_ (
  .A1(_123_),
  .A2(_161_),
  .ZN(_016_)
);

OAI21_X1 _244_ (
  .A(_016_),
  .B1(_123_),
  .B2(_171_),
  .ZN(_017_)
);

NOR2_X1 _245_ (
  .A1(_122_),
  .A2(_017_),
  .ZN(_018_)
);

OAI21_X1 _246_ (
  .A(_011_),
  .B1(_015_),
  .B2(_018_),
  .ZN(_003_)
);

NAND2_X1 _247_ (
  .A1(_116_),
  .A2(\coef[25] ),
  .ZN(_019_)
);

INV_X1 _248_ (
  .A(_163_),
  .ZN(_020_)
);

NAND2_X2 _249_ (
  .A1(_091_),
  .A2(_020_),
  .ZN(_021_)
);

NAND2_X4 _250_ (
  .A1(_123_),
  .A2(_169_),
  .ZN(_022_)
);

NAND3_X2 _251_ (
  .A1(_021_),
  .A2(_103_),
  .A3(_022_),
  .ZN(_023_)
);

NAND2_X2 _252_ (
  .A1(x[0]),
  .A2(_096_),
  .ZN(_024_)
);

NAND2_X1 _253_ (
  .A1(_023_),
  .A2(_024_),
  .ZN(_025_)
);

NAND2_X1 _254_ (
  .A1(_025_),
  .A2(_121_),
  .ZN(_026_)
);

INV_X1 _255_ (
  .A(_165_),
  .ZN(_027_)
);

NAND2_X2 _256_ (
  .A1(_091_),
  .A2(_027_),
  .ZN(_028_)
);

NAND2_X1 _257_ (
  .A1(_090_),
  .A2(_167_),
  .ZN(_029_)
);

NAND3_X1 _258_ (
  .A1(_028_),
  .A2(_097_),
  .A3(_029_),
  .ZN(_030_)
);

INV_X1 _259_ (
  .A(_099_),
  .ZN(_031_)
);

NAND3_X1 _260_ (
  .A1(_030_),
  .A2(_031_),
  .A3(_136_),
  .ZN(_032_)
);

NAND3_X1 _261_ (
  .A1(_026_),
  .A2(_032_),
  .A3(_114_),
  .ZN(_033_)
);

NAND3_X2 _262_ (
  .A1(_021_),
  .A2(_097_),
  .A3(_022_),
  .ZN(_034_)
);

AOI21_X1 _263_ (
  .A(_110_),
  .B1(_034_),
  .B2(_101_),
  .ZN(_035_)
);

NAND2_X2 _264_ (
  .A1(_028_),
  .A2(_029_),
  .ZN(_036_)
);

NAND2_X1 _265_ (
  .A1(_036_),
  .A2(_103_),
  .ZN(_037_)
);

NAND2_X1 _266_ (
  .A1(_037_),
  .A2(_106_),
  .ZN(_038_)
);

AND2_X2 _267_ (
  .A1(_035_),
  .A2(_038_),
  .ZN(_039_)
);

OAI21_X2 _268_ (
  .A(_019_),
  .B1(_033_),
  .B2(_039_),
  .ZN(_004_)
);

NOR2_X1 _269_ (
  .A1(x[0]),
  .A2(_096_),
  .ZN(_040_)
);

NOR2_X1 _270_ (
  .A1(_040_),
  .A2(_120_),
  .ZN(_041_)
);

NAND2_X2 _271_ (
  .A1(_091_),
  .A2(_167_),
  .ZN(_042_)
);

NAND2_X4 _272_ (
  .A1(_027_),
  .A2(_123_),
  .ZN(_043_)
);

NAND2_X4 _273_ (
  .A1(_042_),
  .A2(_043_),
  .ZN(_044_)
);

OAI21_X1 _274_ (
  .A(_041_),
  .B1(_044_),
  .B2(_103_),
  .ZN(_045_)
);

NAND2_X1 _275_ (
  .A1(_024_),
  .A2(_120_),
  .ZN(_046_)
);

INV_X2 _276_ (
  .A(_046_),
  .ZN(_047_)
);

INV_X1 _277_ (
  .A(_169_),
  .ZN(_048_)
);

NAND2_X2 _278_ (
  .A1(_091_),
  .A2(_048_),
  .ZN(_049_)
);

NAND2_X4 _279_ (
  .A1(_123_),
  .A2(_163_),
  .ZN(_050_)
);

NAND2_X4 _280_ (
  .A1(_049_),
  .A2(_050_),
  .ZN(_051_)
);

OAI21_X1 _281_ (
  .A(_047_),
  .B1(_051_),
  .B2(_097_),
  .ZN(_052_)
);

NAND2_X1 _282_ (
  .A1(_045_),
  .A2(_052_),
  .ZN(_053_)
);

NAND2_X1 _283_ (
  .A1(_053_),
  .A2(_109_),
  .ZN(_054_)
);

NAND2_X1 _284_ (
  .A1(_051_),
  .A2(_097_),
  .ZN(_055_)
);

NAND2_X1 _285_ (
  .A1(_055_),
  .A2(_041_),
  .ZN(_056_)
);

NAND2_X1 _286_ (
  .A1(_044_),
  .A2(_103_),
  .ZN(_057_)
);

NAND2_X1 _287_ (
  .A1(_057_),
  .A2(_047_),
  .ZN(_058_)
);

NAND3_X1 _288_ (
  .A1(_056_),
  .A2(_058_),
  .A3(_110_),
  .ZN(_059_)
);

NAND3_X1 _289_ (
  .A1(_054_),
  .A2(_059_),
  .A3(_114_),
  .ZN(_060_)
);

NAND2_X1 _290_ (
  .A1(_116_),
  .A2(\coef[26] ),
  .ZN(_061_)
);

NAND2_X1 _291_ (
  .A1(_060_),
  .A2(_061_),
  .ZN(_005_)
);

NAND2_X1 _292_ (
  .A1(_103_),
  .A2(_158_),
  .ZN(_062_)
);

NAND2_X1 _293_ (
  .A1(_091_),
  .A2(_097_),
  .ZN(_063_)
);

NAND3_X1 _294_ (
  .A1(_062_),
  .A2(_063_),
  .A3(_100_),
  .ZN(_064_)
);

NAND2_X1 _295_ (
  .A1(_103_),
  .A2(_123_),
  .ZN(_065_)
);

NAND2_X1 _296_ (
  .A1(_096_),
  .A2(x[1]),
  .ZN(_066_)
);

NAND3_X1 _297_ (
  .A1(_065_),
  .A2(_066_),
  .A3(_120_),
  .ZN(_067_)
);

NAND2_X1 _298_ (
  .A1(_064_),
  .A2(_067_),
  .ZN(_068_)
);

NAND2_X1 _299_ (
  .A1(_068_),
  .A2(_110_),
  .ZN(_069_)
);

NAND3_X1 _300_ (
  .A1(_064_),
  .A2(_067_),
  .A3(_109_),
  .ZN(_070_)
);

NAND3_X1 _301_ (
  .A1(_069_),
  .A2(_070_),
  .A3(_114_),
  .ZN(_071_)
);

INV_X1 _302_ (
  .A(\coef[27] ),
  .ZN(_072_)
);

OAI21_X1 _303_ (
  .A(_071_),
  .B1(_114_),
  .B2(_072_),
  .ZN(_006_)
);

NOR2_X1 _304_ (
  .A1(_113_),
  .A2(\coef[28] ),
  .ZN(_073_)
);

NAND2_X2 _305_ (
  .A1(_098_),
  .A2(_104_),
  .ZN(_074_)
);

XNOR2_X2 _306_ (
  .A(_074_),
  .B(_109_),
  .ZN(_075_)
);

AOI21_X2 _307_ (
  .A(_073_),
  .B1(_075_),
  .B2(_114_),
  .ZN(_007_)
);

NOR2_X1 _308_ (
  .A1(_113_),
  .A2(\coef[15] ),
  .ZN(_076_)
);

AND2_X1 _309_ (
  .A1(_121_),
  .A2(_024_),
  .ZN(_077_)
);

AOI21_X1 _310_ (
  .A(_116_),
  .B1(_037_),
  .B2(_077_),
  .ZN(_078_)
);

INV_X1 _311_ (
  .A(_040_),
  .ZN(_079_)
);

NAND3_X1 _312_ (
  .A1(_034_),
  .A2(_079_),
  .A3(_136_),
  .ZN(_080_)
);

AND2_X1 _313_ (
  .A1(_078_),
  .A2(_080_),
  .ZN(_081_)
);

NAND2_X1 _314_ (
  .A1(_036_),
  .A2(_097_),
  .ZN(_082_)
);

NAND2_X1 _315_ (
  .A1(_082_),
  .A2(_101_),
  .ZN(_083_)
);

NAND2_X1 _316_ (
  .A1(_023_),
  .A2(_106_),
  .ZN(_084_)
);

NAND2_X1 _317_ (
  .A1(_083_),
  .A2(_084_),
  .ZN(_085_)
);

NAND2_X1 _318_ (
  .A1(_085_),
  .A2(_109_),
  .ZN(_086_)
);

AOI21_X2 _319_ (
  .A(_076_),
  .B1(_081_),
  .B2(_086_),
  .ZN(_008_)
);

NOR2_X1 _320_ (
  .A1(_113_),
  .A2(\coef[30] ),
  .ZN(_087_)
);

NAND2_X1 _321_ (
  .A1(_079_),
  .A2(_024_),
  .ZN(_088_)
);

XNOR2_X1 _322_ (
  .A(_088_),
  .B(_110_),
  .ZN(_089_)
);

AOI21_X1 _323_ (
  .A(_087_),
  .B1(_089_),
  .B2(_114_),
  .ZN(_009_)
);

HA_X1 _324_ (
  .A(_157_),
  .B(_158_),
  .CO(_159_),
  .S(_160_)
);

HA_X1 _325_ (
  .A(_157_),
  .B(_158_),
  .CO(_161_),
  .S(_162_)
);

HA_X1 _326_ (
  .A(_157_),
  .B(x[1]),
  .CO(_163_),
  .S(_164_)
);

HA_X1 _327_ (
  .A(_157_),
  .B(x[1]),
  .CO(_165_),
  .S(_166_)
);

HA_X1 _328_ (
  .A(x[0]),
  .B(_158_),
  .CO(_167_),
  .S(_168_)
);

HA_X1 _329_ (
  .A(x[0]),
  .B(_158_),
  .CO(_169_),
  .S(_170_)
);

HA_X1 _330_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_171_),
  .S(_172_)
);

HA_X1 _331_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_173_),
  .S(_174_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_156_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_155_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_154_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_153_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_152_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_151_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_150_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_149_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_148_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_147_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$94a1b10314722615b96d6c8f661cbb82ecebf320\dctu

module \$paramod$99c498a68fd2923ba65be259bfb6e7d8309d79f4\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _185_ (
  .A(x[1]),
  .ZN(_168_)
);

INV_X1 _186_ (
  .A(x[0]),
  .ZN(_167_)
);

BUF_X2 _187_ (
  .A(y[2]),
  .Z(_098_)
);

INV_X1 _188_ (
  .A(_098_),
  .ZN(_099_)
);

BUF_X2 _189_ (
  .A(_099_),
  .Z(_100_)
);

BUF_X8 _190_ (
  .A(x[2]),
  .Z(_101_)
);

INV_X8 _191_ (
  .A(_101_),
  .ZN(_102_)
);

INV_X1 _192_ (
  .A(_175_),
  .ZN(_103_)
);

NAND2_X2 _193_ (
  .A1(_102_),
  .A2(_103_),
  .ZN(_104_)
);

BUF_X8 _194_ (
  .A(y[0]),
  .Z(_105_)
);

INV_X8 _195_ (
  .A(_105_),
  .ZN(_106_)
);

BUF_X16 _196_ (
  .A(_101_),
  .Z(_107_)
);

NAND2_X4 _197_ (
  .A1(_107_),
  .A2(_177_),
  .ZN(_108_)
);

NAND3_X2 _198_ (
  .A1(_104_),
  .A2(_106_),
  .A3(_108_),
  .ZN(_109_)
);

BUF_X4 _199_ (
  .A(_105_),
  .Z(_110_)
);

NAND2_X1 _200_ (
  .A1(_167_),
  .A2(_110_),
  .ZN(_111_)
);

NAND2_X1 _201_ (
  .A1(_109_),
  .A2(_111_),
  .ZN(_112_)
);

BUF_X2 _202_ (
  .A(y[1]),
  .Z(_113_)
);

BUF_X4 _203_ (
  .A(_113_),
  .Z(_114_)
);

AOI21_X1 _204_ (
  .A(_100_),
  .B1(_112_),
  .B2(_114_),
  .ZN(_115_)
);

INV_X1 _205_ (
  .A(_181_),
  .ZN(_116_)
);

NAND2_X2 _206_ (
  .A1(_102_),
  .A2(_116_),
  .ZN(_117_)
);

NAND2_X1 _207_ (
  .A1(_101_),
  .A2(_171_),
  .ZN(_118_)
);

NAND2_X2 _208_ (
  .A1(_117_),
  .A2(_118_),
  .ZN(_119_)
);

NAND2_X1 _209_ (
  .A1(_119_),
  .A2(_105_),
  .ZN(_120_)
);

OAI21_X1 _210_ (
  .A(_120_),
  .B1(_102_),
  .B2(_110_),
  .ZN(_121_)
);

INV_X2 _211_ (
  .A(_113_),
  .ZN(_122_)
);

NAND2_X1 _212_ (
  .A1(_121_),
  .A2(_122_),
  .ZN(_123_)
);

NAND2_X1 _213_ (
  .A1(_115_),
  .A2(_123_),
  .ZN(_124_)
);

BUF_X2 _214_ (
  .A(ena),
  .Z(_125_)
);

INV_X1 _215_ (
  .A(_183_),
  .ZN(_126_)
);

NAND2_X2 _216_ (
  .A1(_102_),
  .A2(_126_),
  .ZN(_127_)
);

NAND2_X4 _217_ (
  .A1(_107_),
  .A2(_169_),
  .ZN(_128_)
);

NAND2_X2 _218_ (
  .A1(_127_),
  .A2(_128_),
  .ZN(_129_)
);

BUF_X16 _219_ (
  .A(_106_),
  .Z(_130_)
);

NAND2_X1 _220_ (
  .A1(_129_),
  .A2(_130_),
  .ZN(_131_)
);

NAND2_X2 _221_ (
  .A1(_107_),
  .A2(_105_),
  .ZN(_132_)
);

NAND2_X1 _222_ (
  .A1(_132_),
  .A2(_113_),
  .ZN(_133_)
);

INV_X1 _223_ (
  .A(_133_),
  .ZN(_134_)
);

NAND2_X1 _224_ (
  .A1(_131_),
  .A2(_134_),
  .ZN(_135_)
);

INV_X1 _225_ (
  .A(_173_),
  .ZN(_136_)
);

NAND2_X2 _226_ (
  .A1(_102_),
  .A2(_136_),
  .ZN(_137_)
);

NAND2_X1 _227_ (
  .A1(_101_),
  .A2(_179_),
  .ZN(_138_)
);

NAND3_X1 _228_ (
  .A1(_137_),
  .A2(_110_),
  .A3(_138_),
  .ZN(_139_)
);

AOI21_X2 _229_ (
  .A(_113_),
  .B1(_167_),
  .B2(_106_),
  .ZN(_140_)
);

NAND2_X1 _230_ (
  .A1(_139_),
  .A2(_140_),
  .ZN(_141_)
);

NAND3_X1 _231_ (
  .A1(_135_),
  .A2(_141_),
  .A3(_100_),
  .ZN(_142_)
);

NAND3_X1 _232_ (
  .A1(_124_),
  .A2(_125_),
  .A3(_142_),
  .ZN(_143_)
);

INV_X1 _233_ (
  .A(ena),
  .ZN(_144_)
);

NAND2_X1 _234_ (
  .A1(_144_),
  .A2(\coef[21] ),
  .ZN(_145_)
);

NAND2_X1 _235_ (
  .A1(_143_),
  .A2(_145_),
  .ZN(_000_)
);

INV_X1 _236_ (
  .A(_140_),
  .ZN(_146_)
);

NOR2_X1 _237_ (
  .A1(_107_),
  .A2(_110_),
  .ZN(_147_)
);

OAI21_X1 _238_ (
  .A(_146_),
  .B1(_122_),
  .B2(_147_),
  .ZN(_148_)
);

NAND3_X2 _239_ (
  .A1(_104_),
  .A2(_105_),
  .A3(_108_),
  .ZN(_149_)
);

NAND3_X1 _240_ (
  .A1(_148_),
  .A2(_100_),
  .A3(_149_),
  .ZN(_150_)
);

NAND2_X1 _241_ (
  .A1(_105_),
  .A2(x[0]),
  .ZN(_151_)
);

MUX2_X2 _242_ (
  .A(_132_),
  .B(_151_),
  .S(_113_),
  .Z(_152_)
);

NAND2_X1 _243_ (
  .A1(_137_),
  .A2(_138_),
  .ZN(_153_)
);

NAND2_X2 _244_ (
  .A1(_153_),
  .A2(_106_),
  .ZN(_154_)
);

NAND3_X1 _245_ (
  .A1(_152_),
  .A2(_098_),
  .A3(_154_),
  .ZN(_155_)
);

NAND3_X1 _246_ (
  .A1(_150_),
  .A2(_125_),
  .A3(_155_),
  .ZN(_156_)
);

NAND2_X1 _247_ (
  .A1(_144_),
  .A2(\coef[23] ),
  .ZN(_157_)
);

NAND2_X1 _248_ (
  .A1(_156_),
  .A2(_157_),
  .ZN(_001_)
);

XNOR2_X2 _249_ (
  .A(_101_),
  .B(_170_),
  .ZN(_009_)
);

NAND2_X1 _250_ (
  .A1(_009_),
  .A2(_130_),
  .ZN(_010_)
);

NAND2_X1 _251_ (
  .A1(_102_),
  .A2(_110_),
  .ZN(_011_)
);

NAND3_X1 _252_ (
  .A1(_010_),
  .A2(_114_),
  .A3(_011_),
  .ZN(_012_)
);

NAND2_X1 _253_ (
  .A1(_102_),
  .A2(_171_),
  .ZN(_013_)
);

NAND2_X1 _254_ (
  .A1(_116_),
  .A2(_101_),
  .ZN(_014_)
);

NAND2_X1 _255_ (
  .A1(_013_),
  .A2(_014_),
  .ZN(_015_)
);

NAND2_X2 _256_ (
  .A1(_015_),
  .A2(_106_),
  .ZN(_016_)
);

NAND2_X1 _257_ (
  .A1(_016_),
  .A2(_149_),
  .ZN(_017_)
);

NAND2_X1 _258_ (
  .A1(_017_),
  .A2(_122_),
  .ZN(_018_)
);

NAND3_X1 _259_ (
  .A1(_012_),
  .A2(_018_),
  .A3(_100_),
  .ZN(_019_)
);

INV_X1 _260_ (
  .A(_009_),
  .ZN(_020_)
);

NAND2_X2 _261_ (
  .A1(_020_),
  .A2(_110_),
  .ZN(_021_)
);

AOI21_X2 _262_ (
  .A(_113_),
  .B1(_130_),
  .B2(_107_),
  .ZN(_022_)
);

AOI21_X2 _263_ (
  .A(_099_),
  .B1(_021_),
  .B2(_022_),
  .ZN(_023_)
);

INV_X1 _264_ (
  .A(_169_),
  .ZN(_024_)
);

NAND2_X2 _265_ (
  .A1(_102_),
  .A2(_024_),
  .ZN(_025_)
);

NAND2_X4 _266_ (
  .A1(_107_),
  .A2(_183_),
  .ZN(_026_)
);

NAND2_X4 _267_ (
  .A1(_025_),
  .A2(_026_),
  .ZN(_027_)
);

NAND2_X4 _268_ (
  .A1(_027_),
  .A2(_105_),
  .ZN(_028_)
);

NAND2_X1 _269_ (
  .A1(_154_),
  .A2(_028_),
  .ZN(_029_)
);

NAND2_X1 _270_ (
  .A1(_029_),
  .A2(_114_),
  .ZN(_030_)
);

NAND2_X1 _271_ (
  .A1(_023_),
  .A2(_030_),
  .ZN(_031_)
);

NAND3_X1 _272_ (
  .A1(_019_),
  .A2(_031_),
  .A3(_125_),
  .ZN(_032_)
);

NAND2_X1 _273_ (
  .A1(_144_),
  .A2(\coef[24] ),
  .ZN(_033_)
);

NAND2_X1 _274_ (
  .A1(_032_),
  .A2(_033_),
  .ZN(_002_)
);

NAND2_X1 _275_ (
  .A1(_102_),
  .A2(_177_),
  .ZN(_034_)
);

NAND2_X1 _276_ (
  .A1(_103_),
  .A2(_107_),
  .ZN(_035_)
);

NAND3_X1 _277_ (
  .A1(_034_),
  .A2(_035_),
  .A3(_130_),
  .ZN(_036_)
);

NAND3_X1 _278_ (
  .A1(_028_),
  .A2(_036_),
  .A3(_114_),
  .ZN(_037_)
);

NAND3_X1 _279_ (
  .A1(_127_),
  .A2(_105_),
  .A3(_128_),
  .ZN(_038_)
);

NAND3_X1 _280_ (
  .A1(_109_),
  .A2(_038_),
  .A3(_122_),
  .ZN(_039_)
);

NAND2_X1 _281_ (
  .A1(_037_),
  .A2(_039_),
  .ZN(_040_)
);

NAND2_X1 _282_ (
  .A1(_040_),
  .A2(_100_),
  .ZN(_041_)
);

INV_X1 _283_ (
  .A(_179_),
  .ZN(_042_)
);

NAND2_X1 _284_ (
  .A1(_102_),
  .A2(_042_),
  .ZN(_043_)
);

NAND2_X1 _285_ (
  .A1(_107_),
  .A2(_173_),
  .ZN(_044_)
);

NAND3_X1 _286_ (
  .A1(_043_),
  .A2(_105_),
  .A3(_044_),
  .ZN(_045_)
);

NAND2_X1 _287_ (
  .A1(_016_),
  .A2(_045_),
  .ZN(_046_)
);

NAND2_X1 _288_ (
  .A1(_046_),
  .A2(_122_),
  .ZN(_047_)
);

NAND3_X1 _289_ (
  .A1(_117_),
  .A2(_130_),
  .A3(_118_),
  .ZN(_048_)
);

NAND3_X1 _290_ (
  .A1(_139_),
  .A2(_048_),
  .A3(_114_),
  .ZN(_049_)
);

NAND3_X1 _291_ (
  .A1(_047_),
  .A2(_049_),
  .A3(_098_),
  .ZN(_050_)
);

NAND3_X1 _292_ (
  .A1(_041_),
  .A2(_050_),
  .A3(_125_),
  .ZN(_051_)
);

NAND2_X1 _293_ (
  .A1(_144_),
  .A2(\coef[10] ),
  .ZN(_052_)
);

NAND2_X1 _294_ (
  .A1(_051_),
  .A2(_052_),
  .ZN(_003_)
);

OAI21_X1 _295_ (
  .A(_149_),
  .B1(_110_),
  .B2(_129_),
  .ZN(_053_)
);

NAND2_X1 _296_ (
  .A1(_053_),
  .A2(_114_),
  .ZN(_054_)
);

AOI21_X1 _297_ (
  .A(_100_),
  .B1(_140_),
  .B2(_151_),
  .ZN(_055_)
);

NAND2_X1 _298_ (
  .A1(_054_),
  .A2(_055_),
  .ZN(_056_)
);

AOI21_X2 _299_ (
  .A(_122_),
  .B1(_167_),
  .B2(_130_),
  .ZN(_057_)
);

AOI21_X1 _300_ (
  .A(_098_),
  .B1(_057_),
  .B2(_151_),
  .ZN(_058_)
);

NAND2_X1 _301_ (
  .A1(_120_),
  .A2(_154_),
  .ZN(_059_)
);

INV_X1 _302_ (
  .A(_059_),
  .ZN(_060_)
);

OAI21_X1 _303_ (
  .A(_058_),
  .B1(_060_),
  .B2(_114_),
  .ZN(_061_)
);

NAND3_X1 _304_ (
  .A1(_056_),
  .A2(_061_),
  .A3(_125_),
  .ZN(_062_)
);

NAND2_X1 _305_ (
  .A1(_144_),
  .A2(\coef[26] ),
  .ZN(_063_)
);

NAND2_X1 _306_ (
  .A1(_062_),
  .A2(_063_),
  .ZN(_004_)
);

NOR2_X1 _307_ (
  .A1(_125_),
  .A2(\coef[13] ),
  .ZN(_064_)
);

NAND3_X1 _308_ (
  .A1(_021_),
  .A2(_114_),
  .A3(_016_),
  .ZN(_065_)
);

NAND3_X1 _309_ (
  .A1(_034_),
  .A2(_035_),
  .A3(_110_),
  .ZN(_066_)
);

AOI21_X2 _310_ (
  .A(_114_),
  .B1(_130_),
  .B2(x[1]),
  .ZN(_067_)
);

AOI21_X1 _311_ (
  .A(_100_),
  .B1(_066_),
  .B2(_067_),
  .ZN(_068_)
);

AOI21_X1 _312_ (
  .A(_144_),
  .B1(_065_),
  .B2(_068_),
  .ZN(_069_)
);

NAND3_X1 _313_ (
  .A1(_010_),
  .A2(_028_),
  .A3(_122_),
  .ZN(_070_)
);

NAND3_X1 _314_ (
  .A1(_043_),
  .A2(_130_),
  .A3(_044_),
  .ZN(_071_)
);

NAND2_X1 _315_ (
  .A1(_168_),
  .A2(_105_),
  .ZN(_072_)
);

NAND2_X1 _316_ (
  .A1(_072_),
  .A2(_114_),
  .ZN(_073_)
);

INV_X1 _317_ (
  .A(_073_),
  .ZN(_074_)
);

AOI21_X1 _318_ (
  .A(_098_),
  .B1(_071_),
  .B2(_074_),
  .ZN(_075_)
);

NAND2_X1 _319_ (
  .A1(_070_),
  .A2(_075_),
  .ZN(_076_)
);

AOI21_X1 _320_ (
  .A(_064_),
  .B1(_069_),
  .B2(_076_),
  .ZN(_005_)
);

NAND2_X1 _321_ (
  .A1(_067_),
  .A2(_151_),
  .ZN(_077_)
);

NAND3_X1 _322_ (
  .A1(_012_),
  .A2(_100_),
  .A3(_077_),
  .ZN(_078_)
);

NAND2_X1 _323_ (
  .A1(_057_),
  .A2(_072_),
  .ZN(_079_)
);

NAND2_X1 _324_ (
  .A1(_023_),
  .A2(_079_),
  .ZN(_080_)
);

NAND3_X1 _325_ (
  .A1(_078_),
  .A2(_080_),
  .A3(_125_),
  .ZN(_081_)
);

NAND2_X1 _326_ (
  .A1(_144_),
  .A2(\coef[28] ),
  .ZN(_082_)
);

NAND2_X1 _327_ (
  .A1(_081_),
  .A2(_082_),
  .ZN(_006_)
);

OAI21_X2 _328_ (
  .A(_028_),
  .B1(_107_),
  .B2(_110_),
  .ZN(_083_)
);

NAND2_X1 _329_ (
  .A1(_083_),
  .A2(_122_),
  .ZN(_084_)
);

NAND2_X1 _330_ (
  .A1(_129_),
  .A2(_110_),
  .ZN(_085_)
);

AOI21_X1 _331_ (
  .A(_122_),
  .B1(_168_),
  .B2(_130_),
  .ZN(_086_)
);

AOI21_X1 _332_ (
  .A(_100_),
  .B1(_085_),
  .B2(_086_),
  .ZN(_087_)
);

NAND2_X1 _333_ (
  .A1(_084_),
  .A2(_087_),
  .ZN(_088_)
);

NAND2_X1 _334_ (
  .A1(_119_),
  .A2(_130_),
  .ZN(_089_)
);

NAND3_X1 _335_ (
  .A1(_089_),
  .A2(_122_),
  .A3(_072_),
  .ZN(_090_)
);

NAND2_X1 _336_ (
  .A1(_016_),
  .A2(_134_),
  .ZN(_091_)
);

NAND2_X1 _337_ (
  .A1(_090_),
  .A2(_091_),
  .ZN(_092_)
);

NAND2_X1 _338_ (
  .A1(_092_),
  .A2(_100_),
  .ZN(_093_)
);

NAND3_X1 _339_ (
  .A1(_088_),
  .A2(_093_),
  .A3(_125_),
  .ZN(_094_)
);

NAND2_X1 _340_ (
  .A1(_144_),
  .A2(\coef[29] ),
  .ZN(_095_)
);

NAND2_X1 _341_ (
  .A1(_094_),
  .A2(_095_),
  .ZN(_007_)
);

NOR2_X1 _342_ (
  .A1(_125_),
  .A2(\coef[30] ),
  .ZN(_096_)
);

XNOR2_X1 _343_ (
  .A(_107_),
  .B(_098_),
  .ZN(_097_)
);

AOI21_X1 _344_ (
  .A(_096_),
  .B1(_097_),
  .B2(_125_),
  .ZN(_008_)
);

HA_X1 _345_ (
  .A(_167_),
  .B(_168_),
  .CO(_169_),
  .S(_170_)
);

HA_X1 _346_ (
  .A(_167_),
  .B(_168_),
  .CO(_171_),
  .S(_172_)
);

HA_X1 _347_ (
  .A(_167_),
  .B(x[1]),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _348_ (
  .A(_167_),
  .B(x[1]),
  .CO(_175_),
  .S(_176_)
);

HA_X1 _349_ (
  .A(x[0]),
  .B(_168_),
  .CO(_177_),
  .S(_178_)
);

HA_X1 _350_ (
  .A(x[0]),
  .B(_168_),
  .CO(_179_),
  .S(_180_)
);

HA_X1 _351_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_181_),
  .S(_182_)
);

HA_X1 _352_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_183_),
  .S(_184_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_166_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_165_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_164_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_163_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_162_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_161_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_160_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_159_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_158_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$99c498a68fd2923ba65be259bfb6e7d8309d79f4\dctu

module \$paramod$9beaa443332981731011e314e41ebdfa5267d059\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _185_ (
  .A(x[0]),
  .ZN(_167_)
);

INV_X1 _186_ (
  .A(x[1]),
  .ZN(_168_)
);

BUF_X2 _187_ (
  .A(ena),
  .Z(_098_)
);

INV_X2 _188_ (
  .A(_098_),
  .ZN(_099_)
);

CLKBUF_X2 _189_ (
  .A(y[1]),
  .Z(_100_)
);

BUF_X2 _190_ (
  .A(_100_),
  .Z(_101_)
);

BUF_X4 _191_ (
  .A(x[2]),
  .Z(_102_)
);

INV_X8 _192_ (
  .A(_102_),
  .ZN(_103_)
);

NAND2_X2 _193_ (
  .A1(_103_),
  .A2(_170_),
  .ZN(_104_)
);

INV_X1 _194_ (
  .A(_170_),
  .ZN(_105_)
);

BUF_X16 _195_ (
  .A(_102_),
  .Z(_106_)
);

NAND2_X4 _196_ (
  .A1(_105_),
  .A2(_106_),
  .ZN(_107_)
);

NAND2_X4 _197_ (
  .A1(_104_),
  .A2(_107_),
  .ZN(_108_)
);

BUF_X4 _198_ (
  .A(y[0]),
  .Z(_109_)
);

BUF_X4 _199_ (
  .A(_109_),
  .Z(_110_)
);

NOR2_X2 _200_ (
  .A1(_108_),
  .A2(_110_),
  .ZN(_111_)
);

INV_X1 _201_ (
  .A(_179_),
  .ZN(_112_)
);

NAND2_X1 _202_ (
  .A1(_103_),
  .A2(_112_),
  .ZN(_113_)
);

NAND2_X1 _203_ (
  .A1(_106_),
  .A2(_173_),
  .ZN(_114_)
);

NAND3_X1 _204_ (
  .A1(_113_),
  .A2(_110_),
  .A3(_114_),
  .ZN(_115_)
);

INV_X1 _205_ (
  .A(_115_),
  .ZN(_116_)
);

OAI21_X1 _206_ (
  .A(_101_),
  .B1(_111_),
  .B2(_116_),
  .ZN(_117_)
);

NAND2_X1 _207_ (
  .A1(_109_),
  .A2(x[1]),
  .ZN(_118_)
);

INV_X4 _208_ (
  .A(_100_),
  .ZN(_119_)
);

NAND2_X1 _209_ (
  .A1(_118_),
  .A2(_119_),
  .ZN(_120_)
);

INV_X1 _210_ (
  .A(_171_),
  .ZN(_121_)
);

NAND2_X2 _211_ (
  .A1(_103_),
  .A2(_121_),
  .ZN(_122_)
);

NAND2_X4 _212_ (
  .A1(_106_),
  .A2(_181_),
  .ZN(_123_)
);

NAND2_X1 _213_ (
  .A1(_122_),
  .A2(_123_),
  .ZN(_124_)
);

INV_X4 _214_ (
  .A(_109_),
  .ZN(_125_)
);

BUF_X4 _215_ (
  .A(_125_),
  .Z(_126_)
);

AOI21_X1 _216_ (
  .A(_120_),
  .B1(_124_),
  .B2(_126_),
  .ZN(_127_)
);

BUF_X2 _217_ (
  .A(y[2]),
  .Z(_128_)
);

NOR2_X1 _218_ (
  .A1(_127_),
  .A2(_128_),
  .ZN(_129_)
);

AOI21_X1 _219_ (
  .A(_099_),
  .B1(_117_),
  .B2(_129_),
  .ZN(_130_)
);

NAND2_X2 _220_ (
  .A1(_103_),
  .A2(_177_),
  .ZN(_131_)
);

INV_X1 _221_ (
  .A(_175_),
  .ZN(_132_)
);

NAND2_X1 _222_ (
  .A1(_132_),
  .A2(_102_),
  .ZN(_133_)
);

AND2_X2 _223_ (
  .A1(_131_),
  .A2(_133_),
  .ZN(_134_)
);

OR2_X1 _224_ (
  .A1(_134_),
  .A2(_110_),
  .ZN(_135_)
);

BUF_X2 _225_ (
  .A(_119_),
  .Z(_136_)
);

NAND3_X2 _226_ (
  .A1(_104_),
  .A2(_107_),
  .A3(_109_),
  .ZN(_137_)
);

NAND3_X1 _227_ (
  .A1(_135_),
  .A2(_136_),
  .A3(_137_),
  .ZN(_138_)
);

INV_X2 _228_ (
  .A(_128_),
  .ZN(_139_)
);

NAND2_X1 _229_ (
  .A1(_103_),
  .A2(_169_),
  .ZN(_140_)
);

INV_X1 _230_ (
  .A(_183_),
  .ZN(_141_)
);

NAND2_X2 _231_ (
  .A1(_141_),
  .A2(_106_),
  .ZN(_142_)
);

NAND2_X1 _232_ (
  .A1(_140_),
  .A2(_142_),
  .ZN(_143_)
);

NAND2_X1 _233_ (
  .A1(_143_),
  .A2(_110_),
  .ZN(_144_)
);

NOR2_X1 _234_ (
  .A1(_109_),
  .A2(x[1]),
  .ZN(_145_)
);

NOR2_X1 _235_ (
  .A1(_145_),
  .A2(_136_),
  .ZN(_146_)
);

AOI21_X1 _236_ (
  .A(_139_),
  .B1(_144_),
  .B2(_146_),
  .ZN(_147_)
);

NAND2_X1 _237_ (
  .A1(_138_),
  .A2(_147_),
  .ZN(_148_)
);

NAND2_X1 _238_ (
  .A1(_130_),
  .A2(_148_),
  .ZN(_149_)
);

NAND2_X1 _239_ (
  .A1(_099_),
  .A2(\coef[21] ),
  .ZN(_150_)
);

NAND2_X1 _240_ (
  .A1(_149_),
  .A2(_150_),
  .ZN(_000_)
);

NOR2_X1 _241_ (
  .A1(_111_),
  .A2(_128_),
  .ZN(_151_)
);

NAND2_X1 _242_ (
  .A1(_134_),
  .A2(_100_),
  .ZN(_152_)
);

NAND2_X1 _243_ (
  .A1(_152_),
  .A2(_110_),
  .ZN(_153_)
);

NOR2_X1 _244_ (
  .A1(_143_),
  .A2(_101_),
  .ZN(_154_)
);

OAI21_X1 _245_ (
  .A(_151_),
  .B1(_153_),
  .B2(_154_),
  .ZN(_155_)
);

NAND3_X1 _246_ (
  .A1(_122_),
  .A2(_101_),
  .A3(_123_),
  .ZN(_156_)
);

NAND3_X1 _247_ (
  .A1(_113_),
  .A2(_119_),
  .A3(_114_),
  .ZN(_157_)
);

NAND3_X1 _248_ (
  .A1(_156_),
  .A2(_157_),
  .A3(_126_),
  .ZN(_009_)
);

AOI21_X1 _249_ (
  .A(_139_),
  .B1(_108_),
  .B2(_110_),
  .ZN(_010_)
);

NAND2_X1 _250_ (
  .A1(_009_),
  .A2(_010_),
  .ZN(_011_)
);

NAND2_X1 _251_ (
  .A1(_155_),
  .A2(_011_),
  .ZN(_012_)
);

NAND2_X1 _252_ (
  .A1(_012_),
  .A2(_098_),
  .ZN(_013_)
);

NAND2_X1 _253_ (
  .A1(_099_),
  .A2(\coef[23] ),
  .ZN(_014_)
);

NAND2_X1 _254_ (
  .A1(_013_),
  .A2(_014_),
  .ZN(_001_)
);

NAND2_X1 _255_ (
  .A1(_103_),
  .A2(_181_),
  .ZN(_015_)
);

NAND2_X1 _256_ (
  .A1(_121_),
  .A2(_106_),
  .ZN(_016_)
);

NAND3_X1 _257_ (
  .A1(_015_),
  .A2(_016_),
  .A3(_126_),
  .ZN(_017_)
);

NAND3_X2 _258_ (
  .A1(_122_),
  .A2(_109_),
  .A3(_123_),
  .ZN(_018_)
);

NAND2_X1 _259_ (
  .A1(_017_),
  .A2(_018_),
  .ZN(_019_)
);

NAND2_X1 _260_ (
  .A1(_019_),
  .A2(_101_),
  .ZN(_020_)
);

NAND2_X1 _261_ (
  .A1(_125_),
  .A2(x[0]),
  .ZN(_021_)
);

NAND2_X1 _262_ (
  .A1(_137_),
  .A2(_021_),
  .ZN(_022_)
);

NAND2_X1 _263_ (
  .A1(_022_),
  .A2(_136_),
  .ZN(_023_)
);

NAND3_X1 _264_ (
  .A1(_020_),
  .A2(_023_),
  .A3(_128_),
  .ZN(_024_)
);

NAND3_X2 _265_ (
  .A1(_140_),
  .A2(_142_),
  .A3(_126_),
  .ZN(_025_)
);

NAND2_X1 _266_ (
  .A1(_103_),
  .A2(_141_),
  .ZN(_026_)
);

NAND2_X1 _267_ (
  .A1(_106_),
  .A2(_169_),
  .ZN(_027_)
);

NAND3_X1 _268_ (
  .A1(_026_),
  .A2(_110_),
  .A3(_027_),
  .ZN(_028_)
);

NAND3_X2 _269_ (
  .A1(_025_),
  .A2(_028_),
  .A3(_119_),
  .ZN(_029_)
);

NAND2_X2 _270_ (
  .A1(_108_),
  .A2(_126_),
  .ZN(_030_)
);

NAND2_X1 _271_ (
  .A1(_167_),
  .A2(_109_),
  .ZN(_031_)
);

NAND3_X1 _272_ (
  .A1(_030_),
  .A2(_101_),
  .A3(_031_),
  .ZN(_032_)
);

NAND2_X1 _273_ (
  .A1(_029_),
  .A2(_032_),
  .ZN(_033_)
);

NAND2_X1 _274_ (
  .A1(_033_),
  .A2(_139_),
  .ZN(_034_)
);

NAND3_X1 _275_ (
  .A1(_024_),
  .A2(_034_),
  .A3(_098_),
  .ZN(_035_)
);

NAND2_X1 _276_ (
  .A1(_099_),
  .A2(\coef[24] ),
  .ZN(_036_)
);

NAND2_X1 _277_ (
  .A1(_035_),
  .A2(_036_),
  .ZN(_002_)
);

NAND2_X1 _278_ (
  .A1(_168_),
  .A2(_110_),
  .ZN(_037_)
);

NAND3_X2 _279_ (
  .A1(_030_),
  .A2(_136_),
  .A3(_037_),
  .ZN(_038_)
);

INV_X1 _280_ (
  .A(_031_),
  .ZN(_039_)
);

NOR2_X1 _281_ (
  .A1(_106_),
  .A2(_109_),
  .ZN(_040_)
);

OAI21_X1 _282_ (
  .A(_101_),
  .B1(_039_),
  .B2(_040_),
  .ZN(_041_)
);

NAND3_X1 _283_ (
  .A1(_038_),
  .A2(_128_),
  .A3(_041_),
  .ZN(_042_)
);

NAND2_X1 _284_ (
  .A1(_126_),
  .A2(x[1]),
  .ZN(_043_)
);

NAND3_X1 _285_ (
  .A1(_137_),
  .A2(_101_),
  .A3(_043_),
  .ZN(_044_)
);

NAND2_X1 _286_ (
  .A1(_106_),
  .A2(_109_),
  .ZN(_045_)
);

NAND2_X1 _287_ (
  .A1(_021_),
  .A2(_045_),
  .ZN(_046_)
);

NAND2_X1 _288_ (
  .A1(_046_),
  .A2(_136_),
  .ZN(_047_)
);

NAND3_X1 _289_ (
  .A1(_044_),
  .A2(_139_),
  .A3(_047_),
  .ZN(_048_)
);

NAND2_X1 _290_ (
  .A1(_042_),
  .A2(_048_),
  .ZN(_049_)
);

NAND2_X1 _291_ (
  .A1(_049_),
  .A2(_098_),
  .ZN(_050_)
);

NAND2_X1 _292_ (
  .A1(_099_),
  .A2(\coef[10] ),
  .ZN(_051_)
);

NAND2_X1 _293_ (
  .A1(_050_),
  .A2(_051_),
  .ZN(_003_)
);

NAND3_X1 _294_ (
  .A1(_038_),
  .A2(_128_),
  .A3(_152_),
  .ZN(_052_)
);

NAND3_X1 _295_ (
  .A1(_044_),
  .A2(_139_),
  .A3(_157_),
  .ZN(_053_)
);

NAND3_X1 _296_ (
  .A1(_052_),
  .A2(_053_),
  .A3(_098_),
  .ZN(_054_)
);

NAND2_X1 _297_ (
  .A1(_099_),
  .A2(\coef[26] ),
  .ZN(_055_)
);

NAND2_X1 _298_ (
  .A1(_054_),
  .A2(_055_),
  .ZN(_004_)
);

NAND2_X1 _299_ (
  .A1(_099_),
  .A2(\coef[13] ),
  .ZN(_056_)
);

NAND2_X1 _300_ (
  .A1(_112_),
  .A2(_106_),
  .ZN(_057_)
);

NAND2_X1 _301_ (
  .A1(_103_),
  .A2(_173_),
  .ZN(_058_)
);

NAND3_X2 _302_ (
  .A1(_057_),
  .A2(_058_),
  .A3(_126_),
  .ZN(_059_)
);

NAND2_X1 _303_ (
  .A1(_059_),
  .A2(_045_),
  .ZN(_060_)
);

NAND2_X1 _304_ (
  .A1(_060_),
  .A2(_136_),
  .ZN(_061_)
);

NAND2_X1 _305_ (
  .A1(_021_),
  .A2(_100_),
  .ZN(_062_)
);

INV_X1 _306_ (
  .A(_062_),
  .ZN(_063_)
);

AND2_X1 _307_ (
  .A1(_015_),
  .A2(_016_),
  .ZN(_064_)
);

OAI21_X1 _308_ (
  .A(_063_),
  .B1(_064_),
  .B2(_126_),
  .ZN(_065_)
);

NAND3_X1 _309_ (
  .A1(_061_),
  .A2(_065_),
  .A3(_139_),
  .ZN(_066_)
);

NAND2_X1 _310_ (
  .A1(_066_),
  .A2(_098_),
  .ZN(_067_)
);

NAND2_X1 _311_ (
  .A1(_103_),
  .A2(_132_),
  .ZN(_068_)
);

NAND2_X1 _312_ (
  .A1(_106_),
  .A2(_177_),
  .ZN(_069_)
);

NAND3_X1 _313_ (
  .A1(_068_),
  .A2(_109_),
  .A3(_069_),
  .ZN(_070_)
);

INV_X1 _314_ (
  .A(_040_),
  .ZN(_071_)
);

NAND3_X1 _315_ (
  .A1(_070_),
  .A2(_101_),
  .A3(_071_),
  .ZN(_072_)
);

NAND3_X1 _316_ (
  .A1(_026_),
  .A2(_126_),
  .A3(_027_),
  .ZN(_073_)
);

NAND2_X1 _317_ (
  .A1(_110_),
  .A2(x[0]),
  .ZN(_074_)
);

NAND3_X1 _318_ (
  .A1(_073_),
  .A2(_136_),
  .A3(_074_),
  .ZN(_075_)
);

AOI21_X1 _319_ (
  .A(_139_),
  .B1(_072_),
  .B2(_075_),
  .ZN(_076_)
);

OAI21_X2 _320_ (
  .A(_056_),
  .B1(_067_),
  .B2(_076_),
  .ZN(_005_)
);

NAND3_X1 _321_ (
  .A1(_131_),
  .A2(_133_),
  .A3(_110_),
  .ZN(_077_)
);

NAND2_X1 _322_ (
  .A1(_077_),
  .A2(_059_),
  .ZN(_078_)
);

NAND2_X1 _323_ (
  .A1(_078_),
  .A2(_136_),
  .ZN(_079_)
);

NAND3_X1 _324_ (
  .A1(_079_),
  .A2(_020_),
  .A3(_128_),
  .ZN(_080_)
);

NAND3_X1 _325_ (
  .A1(_113_),
  .A2(_126_),
  .A3(_114_),
  .ZN(_081_)
);

NAND3_X1 _326_ (
  .A1(_081_),
  .A2(_070_),
  .A3(_101_),
  .ZN(_082_)
);

NAND2_X1 _327_ (
  .A1(_029_),
  .A2(_082_),
  .ZN(_083_)
);

NAND2_X1 _328_ (
  .A1(_083_),
  .A2(_139_),
  .ZN(_084_)
);

NAND3_X1 _329_ (
  .A1(_080_),
  .A2(_084_),
  .A3(_098_),
  .ZN(_085_)
);

NAND2_X1 _330_ (
  .A1(_099_),
  .A2(\coef[28] ),
  .ZN(_086_)
);

NAND2_X1 _331_ (
  .A1(_085_),
  .A2(_086_),
  .ZN(_006_)
);

NOR2_X1 _332_ (
  .A1(_098_),
  .A2(\coef[29] ),
  .ZN(_087_)
);

NAND2_X1 _333_ (
  .A1(_118_),
  .A2(_101_),
  .ZN(_088_)
);

INV_X1 _334_ (
  .A(_088_),
  .ZN(_089_)
);

AOI21_X1 _335_ (
  .A(_128_),
  .B1(_059_),
  .B2(_089_),
  .ZN(_090_)
);

NAND3_X1 _336_ (
  .A1(_025_),
  .A2(_136_),
  .A3(_031_),
  .ZN(_091_)
);

AOI21_X1 _337_ (
  .A(_099_),
  .B1(_090_),
  .B2(_091_),
  .ZN(_092_)
);

INV_X1 _338_ (
  .A(_145_),
  .ZN(_093_)
);

NAND3_X1 _339_ (
  .A1(_070_),
  .A2(_136_),
  .A3(_093_),
  .ZN(_094_)
);

NAND2_X1 _340_ (
  .A1(_018_),
  .A2(_063_),
  .ZN(_095_)
);

NAND3_X1 _341_ (
  .A1(_094_),
  .A2(_128_),
  .A3(_095_),
  .ZN(_096_)
);

AOI21_X1 _342_ (
  .A(_087_),
  .B1(_092_),
  .B2(_096_),
  .ZN(_007_)
);

NAND2_X1 _343_ (
  .A1(_025_),
  .A2(_018_),
  .ZN(_097_)
);

MUX2_X1 _344_ (
  .A(\coef[30] ),
  .B(_097_),
  .S(_098_),
  .Z(_008_)
);

HA_X1 _345_ (
  .A(_167_),
  .B(_168_),
  .CO(_169_),
  .S(_170_)
);

HA_X1 _346_ (
  .A(_167_),
  .B(_168_),
  .CO(_171_),
  .S(_172_)
);

HA_X1 _347_ (
  .A(_167_),
  .B(x[1]),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _348_ (
  .A(_167_),
  .B(x[1]),
  .CO(_175_),
  .S(_176_)
);

HA_X1 _349_ (
  .A(x[0]),
  .B(_168_),
  .CO(_177_),
  .S(_178_)
);

HA_X1 _350_ (
  .A(x[0]),
  .B(_168_),
  .CO(_179_),
  .S(_180_)
);

HA_X1 _351_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_181_),
  .S(_182_)
);

HA_X1 _352_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_183_),
  .S(_184_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_166_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_165_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_164_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_163_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_162_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_161_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_160_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_159_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_158_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$9beaa443332981731011e314e41ebdfa5267d059\dctu

module \$paramod$9e8342fceac8003655f9e71995b4fdeb8565fbe5\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

BUF_X4 _101_ (
  .A(y[2]),
  .Z(_024_)
);

INV_X1 _102_ (
  .A(x[1]),
  .ZN(_025_)
);

INV_X2 _103_ (
  .A(x[2]),
  .ZN(_026_)
);

NAND2_X2 _104_ (
  .A1(_025_),
  .A2(_026_),
  .ZN(_027_)
);

NAND2_X1 _105_ (
  .A1(x[1]),
  .A2(x[2]),
  .ZN(_028_)
);

NAND2_X2 _106_ (
  .A1(_027_),
  .A2(_028_),
  .ZN(_029_)
);

INV_X2 _107_ (
  .A(y[1]),
  .ZN(_030_)
);

AOI21_X1 _108_ (
  .A(_024_),
  .B1(_029_),
  .B2(_030_),
  .ZN(_031_)
);

BUF_X1 _109_ (
  .A(ena),
  .Z(_032_)
);

CLKBUF_X3 _110_ (
  .A(_032_),
  .Z(_033_)
);

INV_X1 _111_ (
  .A(x[0]),
  .ZN(_034_)
);

NAND2_X4 _112_ (
  .A1(_026_),
  .A2(_034_),
  .ZN(_035_)
);

NAND2_X2 _113_ (
  .A1(x[2]),
  .A2(x[0]),
  .ZN(_036_)
);

NAND2_X4 _114_ (
  .A1(_035_),
  .A2(_036_),
  .ZN(_037_)
);

BUF_X4 _115_ (
  .A(y[1]),
  .Z(_038_)
);

NAND2_X1 _116_ (
  .A1(_037_),
  .A2(_038_),
  .ZN(_039_)
);

NAND3_X1 _117_ (
  .A1(_031_),
  .A2(_033_),
  .A3(_039_),
  .ZN(_040_)
);

INV_X1 _118_ (
  .A(_032_),
  .ZN(_041_)
);

NAND2_X1 _119_ (
  .A1(_041_),
  .A2(\coef[21] ),
  .ZN(_042_)
);

NAND2_X1 _120_ (
  .A1(_024_),
  .A2(_032_),
  .ZN(_043_)
);

NAND2_X2 _121_ (
  .A1(_026_),
  .A2(x[1]),
  .ZN(_044_)
);

NAND2_X1 _122_ (
  .A1(_025_),
  .A2(x[2]),
  .ZN(_045_)
);

NAND2_X4 _123_ (
  .A1(_044_),
  .A2(_045_),
  .ZN(_046_)
);

AOI21_X1 _124_ (
  .A(_043_),
  .B1(_046_),
  .B2(_038_),
  .ZN(_047_)
);

INV_X2 _125_ (
  .A(_037_),
  .ZN(_048_)
);

NAND2_X1 _126_ (
  .A1(_048_),
  .A2(_030_),
  .ZN(_049_)
);

NAND2_X1 _127_ (
  .A1(_047_),
  .A2(_049_),
  .ZN(_050_)
);

NAND3_X1 _128_ (
  .A1(_040_),
  .A2(_042_),
  .A3(_050_),
  .ZN(_000_)
);

BUF_X4 _129_ (
  .A(y[0]),
  .Z(_051_)
);

INV_X2 _130_ (
  .A(_051_),
  .ZN(_052_)
);

NAND2_X4 _131_ (
  .A1(_046_),
  .A2(_052_),
  .ZN(_053_)
);

NAND2_X2 _132_ (
  .A1(_029_),
  .A2(_051_),
  .ZN(_054_)
);

NAND2_X2 _133_ (
  .A1(_053_),
  .A2(_054_),
  .ZN(_055_)
);

MUX2_X2 _134_ (
  .A(\coef[22] ),
  .B(_055_),
  .S(_032_),
  .Z(_001_)
);

NAND3_X1 _135_ (
  .A1(_027_),
  .A2(_051_),
  .A3(_028_),
  .ZN(_056_)
);

NAND3_X2 _136_ (
  .A1(_035_),
  .A2(_052_),
  .A3(_036_),
  .ZN(_057_)
);

NAND2_X2 _137_ (
  .A1(_056_),
  .A2(_057_),
  .ZN(_058_)
);

NAND2_X2 _138_ (
  .A1(_058_),
  .A2(_038_),
  .ZN(_059_)
);

INV_X2 _139_ (
  .A(_024_),
  .ZN(_060_)
);

AOI21_X1 _140_ (
  .A(_060_),
  .B1(_037_),
  .B2(_030_),
  .ZN(_061_)
);

NAND2_X2 _141_ (
  .A1(_059_),
  .A2(_061_),
  .ZN(_062_)
);

NAND3_X1 _142_ (
  .A1(_035_),
  .A2(_051_),
  .A3(_036_),
  .ZN(_063_)
);

NAND3_X2 _143_ (
  .A1(_053_),
  .A2(_063_),
  .A3(_030_),
  .ZN(_064_)
);

AOI21_X4 _144_ (
  .A(_024_),
  .B1(_048_),
  .B2(_038_),
  .ZN(_065_)
);

NAND2_X2 _145_ (
  .A1(_064_),
  .A2(_065_),
  .ZN(_066_)
);

NAND2_X2 _146_ (
  .A1(_062_),
  .A2(_066_),
  .ZN(_067_)
);

NAND2_X2 _147_ (
  .A1(_067_),
  .A2(_033_),
  .ZN(_068_)
);

NAND2_X1 _148_ (
  .A1(_041_),
  .A2(\coef[23] ),
  .ZN(_069_)
);

NAND2_X2 _149_ (
  .A1(_068_),
  .A2(_069_),
  .ZN(_002_)
);

NAND2_X1 _150_ (
  .A1(_041_),
  .A2(\coef[24] ),
  .ZN(_070_)
);

XNOR2_X2 _151_ (
  .A(_060_),
  .B(_038_),
  .ZN(_071_)
);

NAND2_X2 _152_ (
  .A1(_055_),
  .A2(_071_),
  .ZN(_072_)
);

NAND2_X2 _153_ (
  .A1(_072_),
  .A2(_033_),
  .ZN(_073_)
);

OAI21_X1 _154_ (
  .A(_029_),
  .B1(_024_),
  .B2(_038_),
  .ZN(_074_)
);

OAI21_X1 _155_ (
  .A(_046_),
  .B1(_060_),
  .B2(_030_),
  .ZN(_075_)
);

NAND2_X1 _156_ (
  .A1(_074_),
  .A2(_075_),
  .ZN(_076_)
);

INV_X1 _157_ (
  .A(_076_),
  .ZN(_077_)
);

OAI21_X2 _158_ (
  .A(_070_),
  .B1(_073_),
  .B2(_077_),
  .ZN(_003_)
);

AOI21_X1 _159_ (
  .A(_024_),
  .B1(_048_),
  .B2(_030_),
  .ZN(_078_)
);

NAND2_X1 _160_ (
  .A1(_059_),
  .A2(_078_),
  .ZN(_079_)
);

AOI21_X1 _161_ (
  .A(_060_),
  .B1(_037_),
  .B2(_038_),
  .ZN(_080_)
);

NAND2_X1 _162_ (
  .A1(_064_),
  .A2(_080_),
  .ZN(_081_)
);

NAND3_X1 _163_ (
  .A1(_079_),
  .A2(_081_),
  .A3(_033_),
  .ZN(_082_)
);

NAND2_X1 _164_ (
  .A1(_041_),
  .A2(\coef[25] ),
  .ZN(_083_)
);

NAND2_X1 _165_ (
  .A1(_082_),
  .A2(_083_),
  .ZN(_004_)
);

OAI21_X1 _166_ (
  .A(_046_),
  .B1(_051_),
  .B2(_038_),
  .ZN(_084_)
);

NAND3_X1 _167_ (
  .A1(_037_),
  .A2(_052_),
  .A3(_030_),
  .ZN(_085_)
);

NAND3_X1 _168_ (
  .A1(_084_),
  .A2(_085_),
  .A3(_060_),
  .ZN(_086_)
);

OAI21_X1 _169_ (
  .A(_029_),
  .B1(_052_),
  .B2(_030_),
  .ZN(_087_)
);

NAND4_X1 _170_ (
  .A1(_035_),
  .A2(_036_),
  .A3(_051_),
  .A4(_038_),
  .ZN(_088_)
);

NAND3_X1 _171_ (
  .A1(_087_),
  .A2(_088_),
  .A3(_024_),
  .ZN(_089_)
);

NAND2_X1 _172_ (
  .A1(_086_),
  .A2(_089_),
  .ZN(_090_)
);

NAND2_X1 _173_ (
  .A1(_090_),
  .A2(_033_),
  .ZN(_010_)
);

NAND2_X1 _174_ (
  .A1(_041_),
  .A2(\coef[26] ),
  .ZN(_011_)
);

NAND2_X1 _175_ (
  .A1(_010_),
  .A2(_011_),
  .ZN(_005_)
);

NAND2_X1 _176_ (
  .A1(_041_),
  .A2(\coef[27] ),
  .ZN(_012_)
);

NAND2_X1 _177_ (
  .A1(_037_),
  .A2(_051_),
  .ZN(_013_)
);

AOI21_X1 _178_ (
  .A(_071_),
  .B1(_013_),
  .B2(_057_),
  .ZN(_014_)
);

OAI21_X2 _179_ (
  .A(_012_),
  .B1(_073_),
  .B2(_014_),
  .ZN(_006_)
);

NAND3_X1 _180_ (
  .A1(_049_),
  .A2(_033_),
  .A3(_039_),
  .ZN(_015_)
);

INV_X1 _181_ (
  .A(\coef[28] ),
  .ZN(_016_)
);

OAI21_X1 _182_ (
  .A(_015_),
  .B1(_033_),
  .B2(_016_),
  .ZN(_007_)
);

NAND3_X1 _183_ (
  .A1(_053_),
  .A2(_063_),
  .A3(_038_),
  .ZN(_017_)
);

NAND3_X1 _184_ (
  .A1(_017_),
  .A2(_033_),
  .A3(_031_),
  .ZN(_018_)
);

NAND2_X1 _185_ (
  .A1(_058_),
  .A2(_030_),
  .ZN(_019_)
);

NAND2_X1 _186_ (
  .A1(_019_),
  .A2(_047_),
  .ZN(_020_)
);

NAND2_X1 _187_ (
  .A1(_041_),
  .A2(\coef[15] ),
  .ZN(_021_)
);

NAND3_X1 _188_ (
  .A1(_018_),
  .A2(_020_),
  .A3(_021_),
  .ZN(_008_)
);

NOR2_X1 _189_ (
  .A1(_033_),
  .A2(\coef[30] ),
  .ZN(_022_)
);

XNOR2_X1 _190_ (
  .A(_037_),
  .B(_060_),
  .ZN(_023_)
);

AOI21_X1 _191_ (
  .A(_022_),
  .B1(_023_),
  .B2(_033_),
  .ZN(_009_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_100_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_099_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_098_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_097_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_096_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_095_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_094_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_093_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_092_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_091_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$9e8342fceac8003655f9e71995b4fdeb8565fbe5\dctu

module \$paramod$9f831900faf0e9bfdbd9e0f8aa853df59256a109\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _56_ (
  .A(x[0]),
  .ZN(_42_)
);

INV_X1 _57_ (
  .A(x[1]),
  .ZN(_43_)
);

BUF_X4 _58_ (
  .A(ena),
  .Z(_08_)
);

INV_X4 _59_ (
  .A(_08_),
  .ZN(_09_)
);

BUF_X16 _60_ (
  .A(_09_),
  .Z(_10_)
);

NAND2_X4 _61_ (
  .A1(_10_),
  .A2(\coef[21] ),
  .ZN(_11_)
);

BUF_X4 _62_ (
  .A(x[2]),
  .Z(_12_)
);

NAND2_X1 _63_ (
  .A1(_12_),
  .A2(_50_),
  .ZN(_13_)
);

NAND2_X1 _64_ (
  .A1(_13_),
  .A2(_08_),
  .ZN(_14_)
);

NOR2_X1 _65_ (
  .A1(_12_),
  .A2(_48_),
  .ZN(_15_)
);

OAI21_X2 _66_ (
  .A(_11_),
  .B1(_14_),
  .B2(_15_),
  .ZN(_00_)
);

NAND2_X4 _67_ (
  .A1(_10_),
  .A2(\coef[22] ),
  .ZN(_16_)
);

OAI21_X2 _68_ (
  .A(_16_),
  .B1(x[1]),
  .B2(_10_),
  .ZN(_01_)
);

NAND2_X4 _69_ (
  .A1(_10_),
  .A2(\coef[23] ),
  .ZN(_17_)
);

OAI21_X2 _70_ (
  .A(_17_),
  .B1(_12_),
  .B2(_10_),
  .ZN(_02_)
);

NAND2_X4 _71_ (
  .A1(_10_),
  .A2(\coef[14] ),
  .ZN(_18_)
);

OAI21_X2 _72_ (
  .A(_18_),
  .B1(_43_),
  .B2(_10_),
  .ZN(_03_)
);

NAND2_X4 _73_ (
  .A1(_10_),
  .A2(\coef[13] ),
  .ZN(_19_)
);

NAND2_X1 _74_ (
  .A1(_12_),
  .A2(_52_),
  .ZN(_20_)
);

NAND2_X1 _75_ (
  .A1(_20_),
  .A2(_08_),
  .ZN(_21_)
);

NOR2_X1 _76_ (
  .A1(_12_),
  .A2(_46_),
  .ZN(_22_)
);

OAI21_X2 _77_ (
  .A(_19_),
  .B1(_21_),
  .B2(_22_),
  .ZN(_04_)
);

NAND2_X1 _78_ (
  .A1(_09_),
  .A2(\coef[28] ),
  .ZN(_23_)
);

NAND2_X1 _79_ (
  .A1(_12_),
  .A2(_44_),
  .ZN(_24_)
);

NAND2_X1 _80_ (
  .A1(_24_),
  .A2(_08_),
  .ZN(_25_)
);

NOR2_X1 _81_ (
  .A1(_12_),
  .A2(_54_),
  .ZN(_26_)
);

OAI21_X1 _82_ (
  .A(_23_),
  .B1(_25_),
  .B2(_26_),
  .ZN(_05_)
);

INV_X1 _83_ (
  .A(_12_),
  .ZN(_27_)
);

INV_X1 _84_ (
  .A(_45_),
  .ZN(_28_)
);

NAND2_X1 _85_ (
  .A1(_27_),
  .A2(_28_),
  .ZN(_29_)
);

NAND2_X1 _86_ (
  .A1(_12_),
  .A2(_45_),
  .ZN(_30_)
);

NAND3_X1 _87_ (
  .A1(_29_),
  .A2(_08_),
  .A3(_30_),
  .ZN(_31_)
);

NAND2_X4 _88_ (
  .A1(_10_),
  .A2(\coef[15] ),
  .ZN(_32_)
);

NAND2_X2 _89_ (
  .A1(_31_),
  .A2(_32_),
  .ZN(_06_)
);

NAND2_X1 _90_ (
  .A1(_09_),
  .A2(\coef[12] ),
  .ZN(_33_)
);

OAI21_X2 _91_ (
  .A(_33_),
  .B1(_42_),
  .B2(_10_),
  .ZN(_07_)
);

HA_X1 _92_ (
  .A(_42_),
  .B(_43_),
  .CO(_44_),
  .S(_45_)
);

HA_X1 _93_ (
  .A(_42_),
  .B(_43_),
  .CO(_46_),
  .S(_47_)
);

HA_X1 _94_ (
  .A(_42_),
  .B(x[1]),
  .CO(_48_),
  .S(_49_)
);

HA_X1 _95_ (
  .A(x[0]),
  .B(_43_),
  .CO(_50_),
  .S(_51_)
);

HA_X1 _96_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_52_),
  .S(_53_)
);

HA_X1 _97_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_54_),
  .S(_55_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_41_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_01_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_40_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_02_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_39_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_03_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_38_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_04_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_37_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_05_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_36_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_06_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_35_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_07_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_34_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$9f831900faf0e9bfdbd9e0f8aa853df59256a109\dctu

module \$paramod$9fe6c97945bcc341eadabee9cbdea0f75515e5c3\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire \coef[10] ;
wire \coef[11] ;
wire \coef[13] ;
wire \coef[15] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _056_ (
  .A(x[0]),
  .ZN(_004_)
);

BUF_X4 _057_ (
  .A(x[2]),
  .Z(_005_)
);

NAND2_X1 _058_ (
  .A1(_004_),
  .A2(_005_),
  .ZN(_006_)
);

INV_X4 _059_ (
  .A(_005_),
  .ZN(_007_)
);

NAND2_X2 _060_ (
  .A1(_007_),
  .A2(x[0]),
  .ZN(_008_)
);

NAND2_X2 _061_ (
  .A1(_006_),
  .A2(_008_),
  .ZN(_009_)
);

BUF_X4 _062_ (
  .A(y[0]),
  .Z(_010_)
);

INV_X4 _063_ (
  .A(_010_),
  .ZN(_011_)
);

BUF_X4 _064_ (
  .A(y[1]),
  .Z(_012_)
);

INV_X8 _065_ (
  .A(_012_),
  .ZN(_013_)
);

NAND2_X2 _066_ (
  .A1(_011_),
  .A2(_013_),
  .ZN(_014_)
);

NAND2_X1 _067_ (
  .A1(_010_),
  .A2(_012_),
  .ZN(_015_)
);

NAND2_X2 _068_ (
  .A1(_014_),
  .A2(_015_),
  .ZN(_016_)
);

NAND2_X2 _069_ (
  .A1(_009_),
  .A2(_016_),
  .ZN(_017_)
);

NAND2_X2 _070_ (
  .A1(_004_),
  .A2(_007_),
  .ZN(_018_)
);

NAND2_X1 _071_ (
  .A1(x[0]),
  .A2(_005_),
  .ZN(_019_)
);

NAND2_X2 _072_ (
  .A1(_018_),
  .A2(_019_),
  .ZN(_020_)
);

NAND2_X2 _073_ (
  .A1(_011_),
  .A2(_012_),
  .ZN(_021_)
);

NAND2_X2 _074_ (
  .A1(_013_),
  .A2(_010_),
  .ZN(_022_)
);

NAND2_X4 _075_ (
  .A1(_021_),
  .A2(_022_),
  .ZN(_023_)
);

NAND2_X4 _076_ (
  .A1(_020_),
  .A2(_023_),
  .ZN(_024_)
);

CLKBUF_X2 _077_ (
  .A(ena),
  .Z(_025_)
);

NAND3_X1 _078_ (
  .A1(_017_),
  .A2(_024_),
  .A3(_025_),
  .ZN(_026_)
);

INV_X1 _079_ (
  .A(_025_),
  .ZN(_027_)
);

NAND2_X1 _080_ (
  .A1(_027_),
  .A2(\coef[11] ),
  .ZN(_028_)
);

NAND2_X1 _081_ (
  .A1(_026_),
  .A2(_028_),
  .ZN(_000_)
);

INV_X1 _082_ (
  .A(x[1]),
  .ZN(_029_)
);

NAND2_X1 _083_ (
  .A1(_013_),
  .A2(_029_),
  .ZN(_030_)
);

NAND2_X1 _084_ (
  .A1(_012_),
  .A2(x[1]),
  .ZN(_031_)
);

NAND2_X2 _085_ (
  .A1(_030_),
  .A2(_031_),
  .ZN(_032_)
);

NAND2_X1 _086_ (
  .A1(_007_),
  .A2(_010_),
  .ZN(_033_)
);

NAND2_X2 _087_ (
  .A1(_011_),
  .A2(_005_),
  .ZN(_034_)
);

NAND2_X2 _088_ (
  .A1(_033_),
  .A2(_034_),
  .ZN(_035_)
);

NAND2_X4 _089_ (
  .A1(_032_),
  .A2(_035_),
  .ZN(_036_)
);

NAND2_X2 _090_ (
  .A1(_013_),
  .A2(x[1]),
  .ZN(_037_)
);

NAND2_X1 _091_ (
  .A1(_029_),
  .A2(_012_),
  .ZN(_038_)
);

NAND2_X2 _092_ (
  .A1(_037_),
  .A2(_038_),
  .ZN(_039_)
);

NAND2_X2 _093_ (
  .A1(_007_),
  .A2(_011_),
  .ZN(_040_)
);

NAND2_X1 _094_ (
  .A1(_005_),
  .A2(_010_),
  .ZN(_041_)
);

NAND2_X2 _095_ (
  .A1(_040_),
  .A2(_041_),
  .ZN(_042_)
);

NAND2_X4 _096_ (
  .A1(_039_),
  .A2(_042_),
  .ZN(_043_)
);

NAND3_X2 _097_ (
  .A1(_036_),
  .A2(_043_),
  .A3(_025_),
  .ZN(_044_)
);

NAND2_X1 _098_ (
  .A1(_027_),
  .A2(\coef[13] ),
  .ZN(_045_)
);

NAND2_X2 _099_ (
  .A1(_044_),
  .A2(_045_),
  .ZN(_001_)
);

NAND2_X4 _100_ (
  .A1(_036_),
  .A2(_043_),
  .ZN(_046_)
);

NAND2_X4 _101_ (
  .A1(_046_),
  .A2(_025_),
  .ZN(_047_)
);

NAND2_X1 _102_ (
  .A1(_027_),
  .A2(\coef[10] ),
  .ZN(_048_)
);

NAND2_X4 _103_ (
  .A1(_047_),
  .A2(_048_),
  .ZN(_002_)
);

NAND2_X2 _104_ (
  .A1(_017_),
  .A2(_024_),
  .ZN(_049_)
);

NAND2_X2 _105_ (
  .A1(_049_),
  .A2(_025_),
  .ZN(_050_)
);

NAND2_X1 _106_ (
  .A1(_027_),
  .A2(\coef[15] ),
  .ZN(_051_)
);

NAND2_X2 _107_ (
  .A1(_050_),
  .A2(_051_),
  .ZN(_003_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[11] ),
  .QN(_055_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_054_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_053_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_052_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[15] , \coef[15] , \coef[10] , \coef[13] , \coef[10] , \coef[15] , \coef[15] , \coef[11] , \coef[10] , \coef[11] , \coef[15] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$9fe6c97945bcc341eadabee9cbdea0f75515e5c3\dctu

module \$paramod$a184ef4c0e9b8e48eac4b335f6b36fd82c0c32d3\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _095_ (
  .A(x[0]),
  .ZN(_077_)
);

INV_X1 _096_ (
  .A(x[1]),
  .ZN(_078_)
);

BUF_X2 _097_ (
  .A(ena),
  .Z(_012_)
);

NOR2_X1 _098_ (
  .A1(\coef[21] ),
  .A2(_012_),
  .ZN(_013_)
);

INV_X1 _099_ (
  .A(y[0]),
  .ZN(_014_)
);

INV_X1 _100_ (
  .A(y[1]),
  .ZN(_015_)
);

NAND2_X4 _101_ (
  .A1(_014_),
  .A2(_015_),
  .ZN(_016_)
);

NAND2_X1 _102_ (
  .A1(y[0]),
  .A2(y[1]),
  .ZN(_017_)
);

NAND2_X4 _103_ (
  .A1(_016_),
  .A2(_017_),
  .ZN(_018_)
);

XNOR2_X2 _104_ (
  .A(_018_),
  .B(x[1]),
  .ZN(_019_)
);

BUF_X2 _105_ (
  .A(_012_),
  .Z(_020_)
);

AOI21_X1 _106_ (
  .A(_013_),
  .B1(_019_),
  .B2(_020_),
  .ZN(_000_)
);

BUF_X8 _107_ (
  .A(x[2]),
  .Z(_021_)
);

INV_X8 _108_ (
  .A(_021_),
  .ZN(_022_)
);

NAND2_X1 _109_ (
  .A1(_022_),
  .A2(_091_),
  .ZN(_023_)
);

OAI21_X1 _110_ (
  .A(_023_),
  .B1(_022_),
  .B2(_081_),
  .ZN(_024_)
);

NAND2_X1 _111_ (
  .A1(_014_),
  .A2(y[1]),
  .ZN(_025_)
);

NAND2_X1 _112_ (
  .A1(_015_),
  .A2(y[0]),
  .ZN(_026_)
);

NAND2_X2 _113_ (
  .A1(_025_),
  .A2(_026_),
  .ZN(_027_)
);

NAND2_X1 _114_ (
  .A1(_024_),
  .A2(_027_),
  .ZN(_028_)
);

NAND2_X1 _115_ (
  .A1(_021_),
  .A2(_079_),
  .ZN(_029_)
);

OAI21_X1 _116_ (
  .A(_029_),
  .B1(_093_),
  .B2(_021_),
  .ZN(_030_)
);

NAND2_X1 _117_ (
  .A1(_030_),
  .A2(_018_),
  .ZN(_031_)
);

NAND3_X1 _118_ (
  .A1(_028_),
  .A2(_031_),
  .A3(_012_),
  .ZN(_032_)
);

INV_X1 _119_ (
  .A(\coef[22] ),
  .ZN(_033_)
);

OAI21_X1 _120_ (
  .A(_032_),
  .B1(_020_),
  .B2(_033_),
  .ZN(_001_)
);

NAND2_X1 _121_ (
  .A1(_022_),
  .A2(_089_),
  .ZN(_034_)
);

INV_X1 _122_ (
  .A(_083_),
  .ZN(_035_)
);

NAND2_X1 _123_ (
  .A1(_035_),
  .A2(_021_),
  .ZN(_036_)
);

NAND3_X1 _124_ (
  .A1(_027_),
  .A2(_034_),
  .A3(_036_),
  .ZN(_037_)
);

OR2_X1 _125_ (
  .A1(_087_),
  .A2(_021_),
  .ZN(_038_)
);

NAND2_X1 _126_ (
  .A1(_021_),
  .A2(_085_),
  .ZN(_039_)
);

NAND3_X1 _127_ (
  .A1(_018_),
  .A2(_038_),
  .A3(_039_),
  .ZN(_040_)
);

NAND3_X1 _128_ (
  .A1(_037_),
  .A2(_040_),
  .A3(_012_),
  .ZN(_041_)
);

INV_X1 _129_ (
  .A(\coef[23] ),
  .ZN(_042_)
);

OAI21_X1 _130_ (
  .A(_041_),
  .B1(_020_),
  .B2(_042_),
  .ZN(_002_)
);

NAND2_X1 _131_ (
  .A1(_024_),
  .A2(_018_),
  .ZN(_043_)
);

NAND2_X1 _132_ (
  .A1(_030_),
  .A2(_027_),
  .ZN(_044_)
);

NAND3_X1 _133_ (
  .A1(_043_),
  .A2(_044_),
  .A3(_020_),
  .ZN(_045_)
);

INV_X1 _134_ (
  .A(\coef[14] ),
  .ZN(_046_)
);

OAI21_X1 _135_ (
  .A(_045_),
  .B1(_020_),
  .B2(_046_),
  .ZN(_003_)
);

NOR2_X1 _136_ (
  .A1(_012_),
  .A2(\coef[13] ),
  .ZN(_047_)
);

NAND2_X4 _137_ (
  .A1(_018_),
  .A2(_022_),
  .ZN(_048_)
);

NAND3_X1 _138_ (
  .A1(_016_),
  .A2(_021_),
  .A3(_017_),
  .ZN(_049_)
);

NAND2_X2 _139_ (
  .A1(_048_),
  .A2(_049_),
  .ZN(_050_)
);

AOI21_X1 _140_ (
  .A(_047_),
  .B1(_050_),
  .B2(_020_),
  .ZN(_004_)
);

INV_X1 _141_ (
  .A(_080_),
  .ZN(_051_)
);

NAND2_X1 _142_ (
  .A1(_050_),
  .A2(_051_),
  .ZN(_052_)
);

NAND3_X1 _143_ (
  .A1(_048_),
  .A2(_049_),
  .A3(_080_),
  .ZN(_053_)
);

NAND3_X1 _144_ (
  .A1(_052_),
  .A2(_053_),
  .A3(_020_),
  .ZN(_054_)
);

INV_X1 _145_ (
  .A(_012_),
  .ZN(_055_)
);

NAND2_X1 _146_ (
  .A1(_055_),
  .A2(\coef[28] ),
  .ZN(_056_)
);

NAND2_X1 _147_ (
  .A1(_054_),
  .A2(_056_),
  .ZN(_005_)
);

NAND2_X1 _148_ (
  .A1(_022_),
  .A2(_085_),
  .ZN(_057_)
);

OR2_X4 _149_ (
  .A1(_022_),
  .A2(_087_),
  .ZN(_058_)
);

NAND3_X2 _150_ (
  .A1(_027_),
  .A2(_057_),
  .A3(_058_),
  .ZN(_059_)
);

NAND2_X1 _151_ (
  .A1(_022_),
  .A2(_035_),
  .ZN(_060_)
);

NAND2_X1 _152_ (
  .A1(_021_),
  .A2(_089_),
  .ZN(_061_)
);

NAND3_X1 _153_ (
  .A1(_018_),
  .A2(_060_),
  .A3(_061_),
  .ZN(_062_)
);

NAND3_X1 _154_ (
  .A1(_059_),
  .A2(_062_),
  .A3(_020_),
  .ZN(_063_)
);

INV_X1 _155_ (
  .A(\coef[15] ),
  .ZN(_064_)
);

OAI21_X1 _156_ (
  .A(_063_),
  .B1(_020_),
  .B2(_064_),
  .ZN(_006_)
);

NAND2_X1 _157_ (
  .A1(_022_),
  .A2(_081_),
  .ZN(_065_)
);

OR2_X4 _158_ (
  .A1(_022_),
  .A2(_091_),
  .ZN(_066_)
);

NAND3_X2 _159_ (
  .A1(_027_),
  .A2(_065_),
  .A3(_066_),
  .ZN(_067_)
);

OR2_X1 _160_ (
  .A1(_079_),
  .A2(_021_),
  .ZN(_068_)
);

NAND2_X1 _161_ (
  .A1(_093_),
  .A2(_021_),
  .ZN(_008_)
);

NAND3_X1 _162_ (
  .A1(_018_),
  .A2(_068_),
  .A3(_008_),
  .ZN(_009_)
);

NAND3_X1 _163_ (
  .A1(_067_),
  .A2(_009_),
  .A3(_012_),
  .ZN(_010_)
);

INV_X1 _164_ (
  .A(\coef[12] ),
  .ZN(_011_)
);

OAI21_X1 _165_ (
  .A(_010_),
  .B1(_020_),
  .B2(_011_),
  .ZN(_007_)
);

HA_X1 _166_ (
  .A(_077_),
  .B(_078_),
  .CO(_079_),
  .S(_080_)
);

HA_X1 _167_ (
  .A(_077_),
  .B(_078_),
  .CO(_081_),
  .S(_082_)
);

HA_X1 _168_ (
  .A(_077_),
  .B(x[1]),
  .CO(_083_),
  .S(_084_)
);

HA_X1 _169_ (
  .A(_077_),
  .B(x[1]),
  .CO(_085_),
  .S(_086_)
);

HA_X1 _170_ (
  .A(x[0]),
  .B(_078_),
  .CO(_087_),
  .S(_088_)
);

HA_X1 _171_ (
  .A(x[0]),
  .B(_078_),
  .CO(_089_),
  .S(_090_)
);

HA_X1 _172_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_091_),
  .S(_092_)
);

HA_X1 _173_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_093_),
  .S(_094_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_076_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_075_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_074_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_073_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_072_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_071_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_070_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_069_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$a184ef4c0e9b8e48eac4b335f6b36fd82c0c32d3\dctu

module \$paramod$a523c923d4f86f07f4e81f5d8b04b352dfcc17be\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X2 _109_ (
  .A(x[2]),
  .ZN(_032_)
);

INV_X1 _110_ (
  .A(x[0]),
  .ZN(_033_)
);

NAND2_X4 _111_ (
  .A1(_032_),
  .A2(_033_),
  .ZN(_034_)
);

BUF_X4 _112_ (
  .A(y[0]),
  .Z(_035_)
);

INV_X4 _113_ (
  .A(_035_),
  .ZN(_036_)
);

NAND2_X4 _114_ (
  .A1(x[2]),
  .A2(x[0]),
  .ZN(_037_)
);

NAND3_X1 _115_ (
  .A1(_034_),
  .A2(_036_),
  .A3(_037_),
  .ZN(_038_)
);

INV_X1 _116_ (
  .A(x[1]),
  .ZN(_039_)
);

NAND2_X1 _117_ (
  .A1(_032_),
  .A2(_039_),
  .ZN(_040_)
);

NAND2_X1 _118_ (
  .A1(x[2]),
  .A2(x[1]),
  .ZN(_041_)
);

NAND3_X4 _119_ (
  .A1(_040_),
  .A2(_035_),
  .A3(_041_),
  .ZN(_042_)
);

CLKBUF_X3 _120_ (
  .A(y[1]),
  .Z(_043_)
);

NAND3_X1 _121_ (
  .A1(_038_),
  .A2(_042_),
  .A3(_043_),
  .ZN(_044_)
);

NAND2_X4 _122_ (
  .A1(_034_),
  .A2(_037_),
  .ZN(_045_)
);

NAND2_X4 _123_ (
  .A1(_045_),
  .A2(_036_),
  .ZN(_046_)
);

INV_X2 _124_ (
  .A(y[1]),
  .ZN(_047_)
);

NAND3_X1 _125_ (
  .A1(_046_),
  .A2(_042_),
  .A3(_047_),
  .ZN(_048_)
);

BUF_X4 _126_ (
  .A(y[2]),
  .Z(_049_)
);

NAND3_X1 _127_ (
  .A1(_044_),
  .A2(_048_),
  .A3(_049_),
  .ZN(_050_)
);

NAND2_X1 _128_ (
  .A1(_045_),
  .A2(_035_),
  .ZN(_051_)
);

NAND2_X1 _129_ (
  .A1(_039_),
  .A2(x[2]),
  .ZN(_052_)
);

NAND2_X2 _130_ (
  .A1(_032_),
  .A2(x[1]),
  .ZN(_053_)
);

NAND3_X4 _131_ (
  .A1(_052_),
  .A2(_053_),
  .A3(_036_),
  .ZN(_054_)
);

NAND3_X1 _132_ (
  .A1(_051_),
  .A2(_054_),
  .A3(_047_),
  .ZN(_055_)
);

NAND3_X4 _133_ (
  .A1(_034_),
  .A2(_035_),
  .A3(_037_),
  .ZN(_056_)
);

NAND3_X1 _134_ (
  .A1(_054_),
  .A2(_056_),
  .A3(_043_),
  .ZN(_057_)
);

INV_X1 _135_ (
  .A(_049_),
  .ZN(_058_)
);

NAND3_X1 _136_ (
  .A1(_055_),
  .A2(_057_),
  .A3(_058_),
  .ZN(_059_)
);

BUF_X1 _137_ (
  .A(ena),
  .Z(_060_)
);

CLKBUF_X3 _138_ (
  .A(_060_),
  .Z(_061_)
);

NAND3_X1 _139_ (
  .A1(_050_),
  .A2(_059_),
  .A3(_061_),
  .ZN(_062_)
);

INV_X2 _140_ (
  .A(_060_),
  .ZN(_063_)
);

NAND2_X1 _141_ (
  .A1(_063_),
  .A2(\coef[21] ),
  .ZN(_064_)
);

NAND2_X1 _142_ (
  .A1(_062_),
  .A2(_064_),
  .ZN(_000_)
);

NAND2_X1 _143_ (
  .A1(_046_),
  .A2(_056_),
  .ZN(_065_)
);

NAND2_X1 _144_ (
  .A1(_065_),
  .A2(_047_),
  .ZN(_066_)
);

INV_X1 _145_ (
  .A(_045_),
  .ZN(_067_)
);

AOI21_X1 _146_ (
  .A(_049_),
  .B1(_067_),
  .B2(_043_),
  .ZN(_068_)
);

AOI21_X1 _147_ (
  .A(_063_),
  .B1(_066_),
  .B2(_068_),
  .ZN(_069_)
);

NAND2_X1 _148_ (
  .A1(_065_),
  .A2(_043_),
  .ZN(_070_)
);

NAND2_X1 _149_ (
  .A1(_045_),
  .A2(_047_),
  .ZN(_071_)
);

NAND3_X1 _150_ (
  .A1(_070_),
  .A2(_049_),
  .A3(_071_),
  .ZN(_072_)
);

NAND2_X1 _151_ (
  .A1(_069_),
  .A2(_072_),
  .ZN(_073_)
);

NAND2_X1 _152_ (
  .A1(_063_),
  .A2(\coef[22] ),
  .ZN(_074_)
);

NAND2_X1 _153_ (
  .A1(_073_),
  .A2(_074_),
  .ZN(_001_)
);

NAND3_X1 _154_ (
  .A1(_046_),
  .A2(_042_),
  .A3(_043_),
  .ZN(_075_)
);

NAND3_X1 _155_ (
  .A1(_054_),
  .A2(_042_),
  .A3(_047_),
  .ZN(_076_)
);

NAND3_X1 _156_ (
  .A1(_075_),
  .A2(_076_),
  .A3(_049_),
  .ZN(_077_)
);

NAND3_X1 _157_ (
  .A1(_054_),
  .A2(_056_),
  .A3(_047_),
  .ZN(_078_)
);

NAND3_X1 _158_ (
  .A1(_054_),
  .A2(_042_),
  .A3(_043_),
  .ZN(_079_)
);

NAND3_X1 _159_ (
  .A1(_078_),
  .A2(_079_),
  .A3(_058_),
  .ZN(_080_)
);

NAND2_X1 _160_ (
  .A1(_077_),
  .A2(_080_),
  .ZN(_081_)
);

NAND2_X1 _161_ (
  .A1(_081_),
  .A2(_061_),
  .ZN(_082_)
);

NAND2_X1 _162_ (
  .A1(_063_),
  .A2(\coef[23] ),
  .ZN(_083_)
);

NAND2_X1 _163_ (
  .A1(_082_),
  .A2(_083_),
  .ZN(_002_)
);

NAND2_X1 _164_ (
  .A1(_067_),
  .A2(_043_),
  .ZN(_084_)
);

NAND3_X1 _165_ (
  .A1(_084_),
  .A2(_061_),
  .A3(_071_),
  .ZN(_085_)
);

INV_X1 _166_ (
  .A(\coef[24] ),
  .ZN(_086_)
);

OAI21_X1 _167_ (
  .A(_085_),
  .B1(_061_),
  .B2(_086_),
  .ZN(_003_)
);

NAND2_X1 _168_ (
  .A1(_054_),
  .A2(_056_),
  .ZN(_087_)
);

NAND2_X1 _169_ (
  .A1(_087_),
  .A2(_047_),
  .ZN(_088_)
);

NAND3_X1 _170_ (
  .A1(_088_),
  .A2(_079_),
  .A3(_049_),
  .ZN(_089_)
);

NAND3_X1 _171_ (
  .A1(_052_),
  .A2(_053_),
  .A3(_035_),
  .ZN(_090_)
);

NAND3_X1 _172_ (
  .A1(_090_),
  .A2(_038_),
  .A3(_043_),
  .ZN(_091_)
);

NAND3_X1 _173_ (
  .A1(_076_),
  .A2(_091_),
  .A3(_058_),
  .ZN(_092_)
);

NAND3_X1 _174_ (
  .A1(_089_),
  .A2(_092_),
  .A3(_061_),
  .ZN(_093_)
);

NAND2_X1 _175_ (
  .A1(_063_),
  .A2(\coef[25] ),
  .ZN(_094_)
);

NAND2_X1 _176_ (
  .A1(_093_),
  .A2(_094_),
  .ZN(_004_)
);

AOI21_X1 _177_ (
  .A(_063_),
  .B1(_048_),
  .B2(_068_),
  .ZN(_095_)
);

NAND3_X1 _178_ (
  .A1(_057_),
  .A2(_049_),
  .A3(_071_),
  .ZN(_096_)
);

NAND2_X1 _179_ (
  .A1(_095_),
  .A2(_096_),
  .ZN(_097_)
);

INV_X1 _180_ (
  .A(\coef[26] ),
  .ZN(_098_)
);

OAI21_X1 _181_ (
  .A(_097_),
  .B1(_061_),
  .B2(_098_),
  .ZN(_005_)
);

NAND3_X1 _182_ (
  .A1(_051_),
  .A2(_054_),
  .A3(_043_),
  .ZN(_010_)
);

NAND3_X1 _183_ (
  .A1(_010_),
  .A2(_078_),
  .A3(_049_),
  .ZN(_011_)
);

NAND3_X1 _184_ (
  .A1(_038_),
  .A2(_042_),
  .A3(_047_),
  .ZN(_012_)
);

NAND3_X1 _185_ (
  .A1(_075_),
  .A2(_012_),
  .A3(_058_),
  .ZN(_013_)
);

NAND2_X1 _186_ (
  .A1(_011_),
  .A2(_013_),
  .ZN(_014_)
);

NAND2_X1 _187_ (
  .A1(_014_),
  .A2(_061_),
  .ZN(_015_)
);

NAND2_X1 _188_ (
  .A1(_063_),
  .A2(\coef[27] ),
  .ZN(_016_)
);

NAND2_X1 _189_ (
  .A1(_015_),
  .A2(_016_),
  .ZN(_006_)
);

NOR2_X1 _190_ (
  .A1(_060_),
  .A2(\coef[28] ),
  .ZN(_017_)
);

NAND2_X1 _191_ (
  .A1(_058_),
  .A2(_036_),
  .ZN(_018_)
);

NAND2_X1 _192_ (
  .A1(_049_),
  .A2(_035_),
  .ZN(_019_)
);

INV_X1 _193_ (
  .A(_019_),
  .ZN(_020_)
);

OAI21_X1 _194_ (
  .A(_018_),
  .B1(_020_),
  .B2(_043_),
  .ZN(_021_)
);

NAND2_X1 _195_ (
  .A1(_052_),
  .A2(_053_),
  .ZN(_022_)
);

INV_X1 _196_ (
  .A(_022_),
  .ZN(_023_)
);

XNOR2_X1 _197_ (
  .A(_021_),
  .B(_023_),
  .ZN(_024_)
);

AOI21_X1 _198_ (
  .A(_017_),
  .B1(_024_),
  .B2(_061_),
  .ZN(_007_)
);

NAND3_X1 _199_ (
  .A1(_070_),
  .A2(_048_),
  .A3(_049_),
  .ZN(_025_)
);

NAND3_X1 _200_ (
  .A1(_066_),
  .A2(_057_),
  .A3(_058_),
  .ZN(_026_)
);

NAND3_X1 _201_ (
  .A1(_025_),
  .A2(_026_),
  .A3(_061_),
  .ZN(_027_)
);

NAND2_X1 _202_ (
  .A1(_063_),
  .A2(\coef[15] ),
  .ZN(_028_)
);

NAND2_X1 _203_ (
  .A1(_027_),
  .A2(_028_),
  .ZN(_008_)
);

NOR2_X1 _204_ (
  .A1(_060_),
  .A2(\coef[30] ),
  .ZN(_029_)
);

OAI21_X1 _205_ (
  .A(_018_),
  .B1(_020_),
  .B2(_047_),
  .ZN(_030_)
);

XNOR2_X1 _206_ (
  .A(_030_),
  .B(_023_),
  .ZN(_031_)
);

AOI21_X1 _207_ (
  .A(_029_),
  .B1(_031_),
  .B2(_061_),
  .ZN(_009_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_108_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_107_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_106_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_105_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_104_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_103_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_102_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_101_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_100_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_099_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$a523c923d4f86f07f4e81f5d8b04b352dfcc17be\dctu

module \$paramod$a5796bae454a3870edf919a9404bde7ca4192701\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _177_ (
  .A(x[1]),
  .ZN(_160_)
);

INV_X1 _178_ (
  .A(x[0]),
  .ZN(_159_)
);

BUF_X8 _179_ (
  .A(x[2]),
  .Z(_093_)
);

INV_X8 _180_ (
  .A(_093_),
  .ZN(_094_)
);

INV_X2 _181_ (
  .A(y[0]),
  .ZN(_095_)
);

NAND2_X1 _182_ (
  .A1(_094_),
  .A2(_095_),
  .ZN(_096_)
);

NAND2_X1 _183_ (
  .A1(_160_),
  .A2(y[0]),
  .ZN(_097_)
);

INV_X1 _184_ (
  .A(y[1]),
  .ZN(_098_)
);

NAND3_X1 _185_ (
  .A1(_096_),
  .A2(_097_),
  .A3(_098_),
  .ZN(_099_)
);

NAND2_X1 _186_ (
  .A1(_095_),
  .A2(x[1]),
  .ZN(_100_)
);

BUF_X16 _187_ (
  .A(_093_),
  .Z(_101_)
);

BUF_X4 _188_ (
  .A(y[0]),
  .Z(_102_)
);

NAND2_X2 _189_ (
  .A1(_101_),
  .A2(_102_),
  .ZN(_103_)
);

BUF_X4 _190_ (
  .A(y[1]),
  .Z(_104_)
);

NAND3_X1 _191_ (
  .A1(_100_),
  .A2(_103_),
  .A3(_104_),
  .ZN(_105_)
);

NAND2_X1 _192_ (
  .A1(_099_),
  .A2(_105_),
  .ZN(_106_)
);

BUF_X4 _193_ (
  .A(y[2]),
  .Z(_107_)
);

NAND2_X1 _194_ (
  .A1(_106_),
  .A2(_107_),
  .ZN(_108_)
);

INV_X2 _195_ (
  .A(_107_),
  .ZN(_109_)
);

NAND3_X1 _196_ (
  .A1(_099_),
  .A2(_105_),
  .A3(_109_),
  .ZN(_110_)
);

BUF_X1 _197_ (
  .A(ena),
  .Z(_111_)
);

CLKBUF_X3 _198_ (
  .A(_111_),
  .Z(_112_)
);

NAND3_X1 _199_ (
  .A1(_108_),
  .A2(_110_),
  .A3(_112_),
  .ZN(_113_)
);

INV_X1 _200_ (
  .A(\coef[21] ),
  .ZN(_114_)
);

OAI21_X1 _201_ (
  .A(_113_),
  .B1(_114_),
  .B2(_112_),
  .ZN(_000_)
);

NOR2_X1 _202_ (
  .A1(_111_),
  .A2(\coef[22] ),
  .ZN(_115_)
);

NOR2_X2 _203_ (
  .A1(_109_),
  .A2(_104_),
  .ZN(_116_)
);

NOR2_X1 _204_ (
  .A1(_098_),
  .A2(_107_),
  .ZN(_117_)
);

NOR2_X2 _205_ (
  .A1(_116_),
  .A2(_117_),
  .ZN(_118_)
);

XNOR2_X1 _206_ (
  .A(_118_),
  .B(_159_),
  .ZN(_119_)
);

AOI21_X2 _207_ (
  .A(_115_),
  .B1(_119_),
  .B2(_112_),
  .ZN(_001_)
);

NAND2_X1 _208_ (
  .A1(_097_),
  .A2(_104_),
  .ZN(_120_)
);

INV_X1 _209_ (
  .A(_120_),
  .ZN(_121_)
);

NAND2_X1 _210_ (
  .A1(_094_),
  .A2(_171_),
  .ZN(_122_)
);

INV_X1 _211_ (
  .A(_165_),
  .ZN(_123_)
);

NAND2_X1 _212_ (
  .A1(_123_),
  .A2(_093_),
  .ZN(_124_)
);

NAND2_X1 _213_ (
  .A1(_122_),
  .A2(_124_),
  .ZN(_125_)
);

OAI21_X1 _214_ (
  .A(_121_),
  .B1(_125_),
  .B2(_102_),
  .ZN(_126_)
);

BUF_X4 _215_ (
  .A(_095_),
  .Z(_127_)
);

AOI21_X2 _216_ (
  .A(_104_),
  .B1(_127_),
  .B2(x[1]),
  .ZN(_128_)
);

INV_X1 _217_ (
  .A(_169_),
  .ZN(_129_)
);

NAND2_X1 _218_ (
  .A1(_094_),
  .A2(_129_),
  .ZN(_130_)
);

NAND2_X4 _219_ (
  .A1(_101_),
  .A2(_167_),
  .ZN(_131_)
);

NAND2_X2 _220_ (
  .A1(_130_),
  .A2(_131_),
  .ZN(_132_)
);

OAI21_X1 _221_ (
  .A(_128_),
  .B1(_132_),
  .B2(_127_),
  .ZN(_133_)
);

NAND3_X1 _222_ (
  .A1(_126_),
  .A2(_133_),
  .A3(_107_),
  .ZN(_134_)
);

NAND2_X1 _223_ (
  .A1(_132_),
  .A2(_127_),
  .ZN(_135_)
);

NAND2_X1 _224_ (
  .A1(_135_),
  .A2(_121_),
  .ZN(_136_)
);

NAND2_X1 _225_ (
  .A1(_125_),
  .A2(_102_),
  .ZN(_137_)
);

NAND2_X1 _226_ (
  .A1(_137_),
  .A2(_128_),
  .ZN(_138_)
);

NAND2_X1 _227_ (
  .A1(_136_),
  .A2(_138_),
  .ZN(_139_)
);

NAND2_X1 _228_ (
  .A1(_139_),
  .A2(_109_),
  .ZN(_140_)
);

NAND3_X1 _229_ (
  .A1(_134_),
  .A2(_140_),
  .A3(_112_),
  .ZN(_141_)
);

INV_X1 _230_ (
  .A(_111_),
  .ZN(_142_)
);

NAND2_X1 _231_ (
  .A1(_142_),
  .A2(\coef[23] ),
  .ZN(_143_)
);

NAND2_X1 _232_ (
  .A1(_141_),
  .A2(_143_),
  .ZN(_002_)
);

NAND2_X1 _233_ (
  .A1(_142_),
  .A2(\coef[24] ),
  .ZN(_144_)
);

NAND2_X1 _234_ (
  .A1(_129_),
  .A2(_101_),
  .ZN(_145_)
);

NAND2_X1 _235_ (
  .A1(_094_),
  .A2(_167_),
  .ZN(_146_)
);

NAND3_X1 _236_ (
  .A1(_118_),
  .A2(_145_),
  .A3(_146_),
  .ZN(_147_)
);

NAND2_X1 _237_ (
  .A1(_147_),
  .A2(_112_),
  .ZN(_148_)
);

NAND2_X1 _238_ (
  .A1(_101_),
  .A2(_171_),
  .ZN(_010_)
);

OAI21_X1 _239_ (
  .A(_010_),
  .B1(_101_),
  .B2(_165_),
  .ZN(_011_)
);

NOR2_X1 _240_ (
  .A1(_118_),
  .A2(_011_),
  .ZN(_012_)
);

OAI21_X1 _241_ (
  .A(_144_),
  .B1(_148_),
  .B2(_012_),
  .ZN(_003_)
);

NOR2_X1 _242_ (
  .A1(_112_),
  .A2(\coef[25] ),
  .ZN(_013_)
);

NAND2_X1 _243_ (
  .A1(_094_),
  .A2(_173_),
  .ZN(_014_)
);

INV_X1 _244_ (
  .A(_163_),
  .ZN(_015_)
);

NAND2_X2 _245_ (
  .A1(_015_),
  .A2(_101_),
  .ZN(_016_)
);

NAND3_X2 _246_ (
  .A1(_014_),
  .A2(_016_),
  .A3(_127_),
  .ZN(_017_)
);

NAND2_X1 _247_ (
  .A1(_017_),
  .A2(_103_),
  .ZN(_018_)
);

NAND2_X1 _248_ (
  .A1(_104_),
  .A2(_107_),
  .ZN(_019_)
);

INV_X1 _249_ (
  .A(_019_),
  .ZN(_020_)
);

NAND2_X1 _250_ (
  .A1(_018_),
  .A2(_020_),
  .ZN(_021_)
);

INV_X1 _251_ (
  .A(_175_),
  .ZN(_022_)
);

NAND2_X1 _252_ (
  .A1(_094_),
  .A2(_022_),
  .ZN(_023_)
);

NAND2_X1 _253_ (
  .A1(_093_),
  .A2(_161_),
  .ZN(_024_)
);

NAND3_X2 _254_ (
  .A1(_023_),
  .A2(_127_),
  .A3(_024_),
  .ZN(_025_)
);

NAND2_X1 _255_ (
  .A1(_094_),
  .A2(_102_),
  .ZN(_026_)
);

NAND2_X1 _256_ (
  .A1(_025_),
  .A2(_026_),
  .ZN(_027_)
);

NAND2_X1 _257_ (
  .A1(_027_),
  .A2(_117_),
  .ZN(_028_)
);

NAND2_X1 _258_ (
  .A1(_021_),
  .A2(_028_),
  .ZN(_029_)
);

INV_X1 _259_ (
  .A(_116_),
  .ZN(_030_)
);

NAND3_X1 _260_ (
  .A1(_023_),
  .A2(_102_),
  .A3(_024_),
  .ZN(_031_)
);

AOI21_X1 _261_ (
  .A(_030_),
  .B1(_031_),
  .B2(_096_),
  .ZN(_032_)
);

NOR2_X2 _262_ (
  .A1(_029_),
  .A2(_032_),
  .ZN(_033_)
);

NAND3_X1 _263_ (
  .A1(_014_),
  .A2(_016_),
  .A3(_102_),
  .ZN(_034_)
);

NAND2_X1 _264_ (
  .A1(_095_),
  .A2(_101_),
  .ZN(_035_)
);

NAND2_X1 _265_ (
  .A1(_034_),
  .A2(_035_),
  .ZN(_036_)
);

NOR2_X1 _266_ (
  .A1(_104_),
  .A2(_107_),
  .ZN(_037_)
);

AOI21_X1 _267_ (
  .A(_142_),
  .B1(_036_),
  .B2(_037_),
  .ZN(_038_)
);

AOI21_X2 _268_ (
  .A(_013_),
  .B1(_033_),
  .B2(_038_),
  .ZN(_004_)
);

OR2_X4 _269_ (
  .A1(_161_),
  .A2(_101_),
  .ZN(_039_)
);

NAND2_X1 _270_ (
  .A1(_101_),
  .A2(_175_),
  .ZN(_040_)
);

NAND3_X1 _271_ (
  .A1(_039_),
  .A2(_127_),
  .A3(_040_),
  .ZN(_041_)
);

NAND2_X1 _272_ (
  .A1(_103_),
  .A2(_098_),
  .ZN(_042_)
);

INV_X1 _273_ (
  .A(_042_),
  .ZN(_043_)
);

NAND2_X1 _274_ (
  .A1(_041_),
  .A2(_043_),
  .ZN(_044_)
);

NAND2_X1 _275_ (
  .A1(_094_),
  .A2(_163_),
  .ZN(_045_)
);

INV_X1 _276_ (
  .A(_173_),
  .ZN(_046_)
);

NAND2_X1 _277_ (
  .A1(_046_),
  .A2(_101_),
  .ZN(_047_)
);

NAND3_X1 _278_ (
  .A1(_045_),
  .A2(_047_),
  .A3(_102_),
  .ZN(_048_)
);

AOI21_X1 _279_ (
  .A(_098_),
  .B1(_127_),
  .B2(_094_),
  .ZN(_049_)
);

NAND2_X1 _280_ (
  .A1(_048_),
  .A2(_049_),
  .ZN(_050_)
);

NAND3_X1 _281_ (
  .A1(_044_),
  .A2(_050_),
  .A3(_109_),
  .ZN(_051_)
);

NAND3_X2 _282_ (
  .A1(_039_),
  .A2(_102_),
  .A3(_040_),
  .ZN(_052_)
);

NAND2_X1 _283_ (
  .A1(_035_),
  .A2(_104_),
  .ZN(_053_)
);

INV_X1 _284_ (
  .A(_053_),
  .ZN(_054_)
);

NAND2_X1 _285_ (
  .A1(_052_),
  .A2(_054_),
  .ZN(_055_)
);

NAND3_X1 _286_ (
  .A1(_045_),
  .A2(_047_),
  .A3(_127_),
  .ZN(_056_)
);

AOI21_X1 _287_ (
  .A(_104_),
  .B1(_094_),
  .B2(_102_),
  .ZN(_057_)
);

NAND2_X1 _288_ (
  .A1(_056_),
  .A2(_057_),
  .ZN(_058_)
);

NAND3_X1 _289_ (
  .A1(_055_),
  .A2(_058_),
  .A3(_107_),
  .ZN(_059_)
);

NAND3_X1 _290_ (
  .A1(_051_),
  .A2(_059_),
  .A3(_112_),
  .ZN(_060_)
);

NAND2_X1 _291_ (
  .A1(_142_),
  .A2(\coef[26] ),
  .ZN(_061_)
);

NAND2_X1 _292_ (
  .A1(_060_),
  .A2(_061_),
  .ZN(_005_)
);

OR2_X4 _293_ (
  .A1(_162_),
  .A2(_093_),
  .ZN(_062_)
);

NAND2_X1 _294_ (
  .A1(_093_),
  .A2(_162_),
  .ZN(_063_)
);

NAND2_X2 _295_ (
  .A1(_062_),
  .A2(_063_),
  .ZN(_064_)
);

NAND2_X1 _296_ (
  .A1(_064_),
  .A2(_127_),
  .ZN(_065_)
);

OAI21_X1 _297_ (
  .A(_104_),
  .B1(_095_),
  .B2(_159_),
  .ZN(_066_)
);

INV_X1 _298_ (
  .A(_066_),
  .ZN(_067_)
);

NAND2_X2 _299_ (
  .A1(_065_),
  .A2(_067_),
  .ZN(_068_)
);

NAND3_X1 _300_ (
  .A1(_062_),
  .A2(_102_),
  .A3(_063_),
  .ZN(_069_)
);

AOI21_X2 _301_ (
  .A(_104_),
  .B1(_159_),
  .B2(_127_),
  .ZN(_070_)
);

NAND2_X1 _302_ (
  .A1(_069_),
  .A2(_070_),
  .ZN(_071_)
);

NAND2_X1 _303_ (
  .A1(_068_),
  .A2(_071_),
  .ZN(_072_)
);

NAND2_X1 _304_ (
  .A1(_072_),
  .A2(_109_),
  .ZN(_073_)
);

NAND3_X1 _305_ (
  .A1(_068_),
  .A2(_071_),
  .A3(_107_),
  .ZN(_074_)
);

NAND3_X1 _306_ (
  .A1(_073_),
  .A2(_074_),
  .A3(_112_),
  .ZN(_075_)
);

NAND2_X1 _307_ (
  .A1(_142_),
  .A2(\coef[27] ),
  .ZN(_076_)
);

NAND2_X1 _308_ (
  .A1(_075_),
  .A2(_076_),
  .ZN(_006_)
);

NOR2_X1 _309_ (
  .A1(_111_),
  .A2(\coef[28] ),
  .ZN(_077_)
);

NAND2_X1 _310_ (
  .A1(_100_),
  .A2(_097_),
  .ZN(_078_)
);

XNOR2_X1 _311_ (
  .A(_078_),
  .B(_109_),
  .ZN(_079_)
);

AOI21_X1 _312_ (
  .A(_077_),
  .B1(_079_),
  .B2(_112_),
  .ZN(_007_)
);

NOR2_X1 _313_ (
  .A1(_111_),
  .A2(\coef[15] ),
  .ZN(_080_)
);

NAND2_X1 _314_ (
  .A1(_017_),
  .A2(_026_),
  .ZN(_081_)
);

NAND2_X1 _315_ (
  .A1(_081_),
  .A2(_117_),
  .ZN(_082_)
);

NAND2_X1 _316_ (
  .A1(_025_),
  .A2(_103_),
  .ZN(_083_)
);

NAND2_X1 _317_ (
  .A1(_083_),
  .A2(_020_),
  .ZN(_084_)
);

NAND2_X1 _318_ (
  .A1(_082_),
  .A2(_084_),
  .ZN(_085_)
);

AOI21_X1 _319_ (
  .A(_030_),
  .B1(_034_),
  .B2(_096_),
  .ZN(_086_)
);

NOR2_X2 _320_ (
  .A1(_085_),
  .A2(_086_),
  .ZN(_087_)
);

NAND2_X1 _321_ (
  .A1(_031_),
  .A2(_035_),
  .ZN(_088_)
);

AOI21_X1 _322_ (
  .A(_142_),
  .B1(_088_),
  .B2(_037_),
  .ZN(_089_)
);

AOI21_X2 _323_ (
  .A(_080_),
  .B1(_087_),
  .B2(_089_),
  .ZN(_008_)
);

NOR2_X1 _324_ (
  .A1(_111_),
  .A2(\coef[30] ),
  .ZN(_090_)
);

NAND2_X1 _325_ (
  .A1(_096_),
  .A2(_103_),
  .ZN(_091_)
);

XNOR2_X1 _326_ (
  .A(_091_),
  .B(_109_),
  .ZN(_092_)
);

AOI21_X1 _327_ (
  .A(_090_),
  .B1(_092_),
  .B2(_112_),
  .ZN(_009_)
);

HA_X1 _328_ (
  .A(_159_),
  .B(_160_),
  .CO(_161_),
  .S(_162_)
);

HA_X1 _329_ (
  .A(_159_),
  .B(_160_),
  .CO(_163_),
  .S(_164_)
);

HA_X1 _330_ (
  .A(_159_),
  .B(x[1]),
  .CO(_165_),
  .S(_166_)
);

HA_X1 _331_ (
  .A(_159_),
  .B(x[1]),
  .CO(_167_),
  .S(_168_)
);

HA_X1 _332_ (
  .A(x[0]),
  .B(_160_),
  .CO(_169_),
  .S(_170_)
);

HA_X1 _333_ (
  .A(x[0]),
  .B(_160_),
  .CO(_171_),
  .S(_172_)
);

HA_X1 _334_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _335_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_175_),
  .S(_176_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_158_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_157_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_156_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_155_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_154_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_153_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_152_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_151_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_150_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_149_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$a5796bae454a3870edf919a9404bde7ca4192701\dctu

module \$paramod$a8d3b7b4edaf7d596a54a187c8ed4a9561fa625a\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

BUF_X4 _118_ (
  .A(x[2]),
  .Z(_041_)
);

INV_X8 _119_ (
  .A(_041_),
  .ZN(_042_)
);

NAND2_X4 _120_ (
  .A1(_042_),
  .A2(x[1]),
  .ZN(_043_)
);

INV_X2 _121_ (
  .A(x[1]),
  .ZN(_044_)
);

NAND2_X2 _122_ (
  .A1(_044_),
  .A2(_041_),
  .ZN(_045_)
);

NAND2_X4 _123_ (
  .A1(_043_),
  .A2(_045_),
  .ZN(_046_)
);

NAND2_X4 _124_ (
  .A1(_046_),
  .A2(y[0]),
  .ZN(_047_)
);

INV_X2 _125_ (
  .A(x[0]),
  .ZN(_048_)
);

NAND2_X2 _126_ (
  .A1(_048_),
  .A2(_041_),
  .ZN(_049_)
);

NAND2_X4 _127_ (
  .A1(_042_),
  .A2(x[0]),
  .ZN(_050_)
);

INV_X2 _128_ (
  .A(y[0]),
  .ZN(_051_)
);

NAND3_X2 _129_ (
  .A1(_049_),
  .A2(_050_),
  .A3(_051_),
  .ZN(_052_)
);

BUF_X4 _130_ (
  .A(y[1]),
  .Z(_053_)
);

NAND3_X1 _131_ (
  .A1(_047_),
  .A2(_052_),
  .A3(_053_),
  .ZN(_054_)
);

NAND2_X4 _132_ (
  .A1(_048_),
  .A2(_042_),
  .ZN(_055_)
);

NAND2_X2 _133_ (
  .A1(x[0]),
  .A2(_041_),
  .ZN(_056_)
);

NAND3_X2 _134_ (
  .A1(_055_),
  .A2(_051_),
  .A3(_056_),
  .ZN(_057_)
);

INV_X2 _135_ (
  .A(_053_),
  .ZN(_058_)
);

NAND3_X2 _136_ (
  .A1(_047_),
  .A2(_057_),
  .A3(_058_),
  .ZN(_059_)
);

NAND2_X1 _137_ (
  .A1(_054_),
  .A2(_059_),
  .ZN(_060_)
);

BUF_X2 _138_ (
  .A(y[2]),
  .Z(_061_)
);

INV_X2 _139_ (
  .A(_061_),
  .ZN(_062_)
);

NAND2_X1 _140_ (
  .A1(_060_),
  .A2(_062_),
  .ZN(_063_)
);

NAND3_X2 _141_ (
  .A1(_049_),
  .A2(_050_),
  .A3(y[0]),
  .ZN(_064_)
);

NAND2_X4 _142_ (
  .A1(_042_),
  .A2(_044_),
  .ZN(_065_)
);

NAND2_X1 _143_ (
  .A1(_041_),
  .A2(x[1]),
  .ZN(_066_)
);

NAND3_X1 _144_ (
  .A1(_065_),
  .A2(_051_),
  .A3(_066_),
  .ZN(_067_)
);

BUF_X4 _145_ (
  .A(_058_),
  .Z(_068_)
);

NAND3_X1 _146_ (
  .A1(_064_),
  .A2(_067_),
  .A3(_068_),
  .ZN(_069_)
);

NAND3_X2 _147_ (
  .A1(_055_),
  .A2(y[0]),
  .A3(_056_),
  .ZN(_070_)
);

NAND3_X2 _148_ (
  .A1(_070_),
  .A2(_067_),
  .A3(_053_),
  .ZN(_071_)
);

NAND3_X1 _149_ (
  .A1(_069_),
  .A2(_071_),
  .A3(_061_),
  .ZN(_072_)
);

NAND2_X1 _150_ (
  .A1(_063_),
  .A2(_072_),
  .ZN(_073_)
);

CLKBUF_X3 _151_ (
  .A(ena),
  .Z(_074_)
);

NAND2_X1 _152_ (
  .A1(_073_),
  .A2(_074_),
  .ZN(_075_)
);

INV_X1 _153_ (
  .A(ena),
  .ZN(_076_)
);

NAND2_X1 _154_ (
  .A1(_076_),
  .A2(\coef[21] ),
  .ZN(_077_)
);

NAND2_X2 _155_ (
  .A1(_075_),
  .A2(_077_),
  .ZN(_000_)
);

NAND2_X1 _156_ (
  .A1(_076_),
  .A2(\coef[22] ),
  .ZN(_078_)
);

NAND3_X2 _157_ (
  .A1(_064_),
  .A2(_057_),
  .A3(_053_),
  .ZN(_079_)
);

NAND2_X1 _158_ (
  .A1(_049_),
  .A2(_050_),
  .ZN(_080_)
);

NAND2_X1 _159_ (
  .A1(_080_),
  .A2(_068_),
  .ZN(_081_)
);

AOI21_X1 _160_ (
  .A(_062_),
  .B1(_079_),
  .B2(_081_),
  .ZN(_082_)
);

NAND3_X2 _161_ (
  .A1(_052_),
  .A2(_070_),
  .A3(_058_),
  .ZN(_083_)
);

AOI21_X1 _162_ (
  .A(_061_),
  .B1(_080_),
  .B2(_053_),
  .ZN(_084_)
);

NAND2_X1 _163_ (
  .A1(_083_),
  .A2(_084_),
  .ZN(_085_)
);

NAND2_X1 _164_ (
  .A1(_085_),
  .A2(_074_),
  .ZN(_086_)
);

OAI21_X1 _165_ (
  .A(_078_),
  .B1(_082_),
  .B2(_086_),
  .ZN(_001_)
);

NOR2_X1 _166_ (
  .A1(_074_),
  .A2(\coef[23] ),
  .ZN(_087_)
);

NAND2_X2 _167_ (
  .A1(_065_),
  .A2(_066_),
  .ZN(_088_)
);

NAND2_X2 _168_ (
  .A1(_088_),
  .A2(_051_),
  .ZN(_089_)
);

NAND3_X1 _169_ (
  .A1(_089_),
  .A2(_064_),
  .A3(_068_),
  .ZN(_090_)
);

AOI21_X1 _170_ (
  .A(_062_),
  .B1(_046_),
  .B2(_053_),
  .ZN(_091_)
);

AOI21_X1 _171_ (
  .A(_076_),
  .B1(_090_),
  .B2(_091_),
  .ZN(_092_)
);

NAND3_X1 _172_ (
  .A1(_047_),
  .A2(_057_),
  .A3(_053_),
  .ZN(_093_)
);

AOI21_X1 _173_ (
  .A(_061_),
  .B1(_088_),
  .B2(_068_),
  .ZN(_094_)
);

NAND2_X1 _174_ (
  .A1(_093_),
  .A2(_094_),
  .ZN(_095_)
);

AOI21_X1 _175_ (
  .A(_087_),
  .B1(_092_),
  .B2(_095_),
  .ZN(_002_)
);

NAND2_X1 _176_ (
  .A1(_079_),
  .A2(_083_),
  .ZN(_096_)
);

NAND2_X1 _177_ (
  .A1(_096_),
  .A2(_062_),
  .ZN(_097_)
);

NAND3_X1 _178_ (
  .A1(_079_),
  .A2(_083_),
  .A3(_061_),
  .ZN(_098_)
);

NAND3_X1 _179_ (
  .A1(_097_),
  .A2(_098_),
  .A3(_074_),
  .ZN(_099_)
);

NAND2_X1 _180_ (
  .A1(_076_),
  .A2(\coef[24] ),
  .ZN(_100_)
);

NAND2_X1 _181_ (
  .A1(_099_),
  .A2(_100_),
  .ZN(_003_)
);

NOR2_X1 _182_ (
  .A1(_046_),
  .A2(_068_),
  .ZN(_101_)
);

INV_X1 _183_ (
  .A(_101_),
  .ZN(_102_)
);

NAND3_X1 _184_ (
  .A1(_090_),
  .A2(_062_),
  .A3(_102_),
  .ZN(_103_)
);

NAND2_X1 _185_ (
  .A1(_046_),
  .A2(_068_),
  .ZN(_104_)
);

NAND3_X1 _186_ (
  .A1(_093_),
  .A2(_061_),
  .A3(_104_),
  .ZN(_105_)
);

NAND3_X1 _187_ (
  .A1(_103_),
  .A2(_105_),
  .A3(_074_),
  .ZN(_106_)
);

NAND2_X1 _188_ (
  .A1(_076_),
  .A2(\coef[25] ),
  .ZN(_107_)
);

NAND2_X1 _189_ (
  .A1(_106_),
  .A2(_107_),
  .ZN(_004_)
);

NAND2_X1 _190_ (
  .A1(_071_),
  .A2(_083_),
  .ZN(_010_)
);

NAND2_X1 _191_ (
  .A1(_010_),
  .A2(_062_),
  .ZN(_011_)
);

NAND3_X1 _192_ (
  .A1(_059_),
  .A2(_079_),
  .A3(_061_),
  .ZN(_012_)
);

NAND2_X1 _193_ (
  .A1(_011_),
  .A2(_012_),
  .ZN(_013_)
);

NAND2_X1 _194_ (
  .A1(_013_),
  .A2(_074_),
  .ZN(_014_)
);

NAND2_X1 _195_ (
  .A1(_076_),
  .A2(\coef[26] ),
  .ZN(_015_)
);

NAND2_X1 _196_ (
  .A1(_014_),
  .A2(_015_),
  .ZN(_005_)
);

NAND3_X1 _197_ (
  .A1(_047_),
  .A2(_052_),
  .A3(_068_),
  .ZN(_016_)
);

NAND3_X1 _198_ (
  .A1(_016_),
  .A2(_093_),
  .A3(_061_),
  .ZN(_017_)
);

NAND3_X1 _199_ (
  .A1(_089_),
  .A2(_070_),
  .A3(_053_),
  .ZN(_018_)
);

NAND3_X1 _200_ (
  .A1(_090_),
  .A2(_018_),
  .A3(_062_),
  .ZN(_019_)
);

NAND3_X1 _201_ (
  .A1(_017_),
  .A2(_019_),
  .A3(_074_),
  .ZN(_020_)
);

NAND2_X1 _202_ (
  .A1(_076_),
  .A2(\coef[27] ),
  .ZN(_021_)
);

NAND2_X1 _203_ (
  .A1(_020_),
  .A2(_021_),
  .ZN(_006_)
);

AND2_X4 _204_ (
  .A1(_047_),
  .A2(_089_),
  .ZN(_022_)
);

NAND2_X1 _205_ (
  .A1(_022_),
  .A2(_053_),
  .ZN(_023_)
);

NAND2_X1 _206_ (
  .A1(_023_),
  .A2(_094_),
  .ZN(_024_)
);

NAND2_X1 _207_ (
  .A1(_022_),
  .A2(_068_),
  .ZN(_025_)
);

NAND2_X1 _208_ (
  .A1(_025_),
  .A2(_091_),
  .ZN(_026_)
);

NAND3_X1 _209_ (
  .A1(_024_),
  .A2(_026_),
  .A3(_074_),
  .ZN(_027_)
);

NAND2_X1 _210_ (
  .A1(_076_),
  .A2(\coef[28] ),
  .ZN(_028_)
);

NAND2_X1 _211_ (
  .A1(_027_),
  .A2(_028_),
  .ZN(_007_)
);

NOR2_X1 _212_ (
  .A1(_074_),
  .A2(\coef[15] ),
  .ZN(_029_)
);

AOI21_X1 _213_ (
  .A(_062_),
  .B1(_080_),
  .B2(_068_),
  .ZN(_030_)
);

AOI21_X1 _214_ (
  .A(_076_),
  .B1(_071_),
  .B2(_030_),
  .ZN(_031_)
);

NAND2_X1 _215_ (
  .A1(_080_),
  .A2(_053_),
  .ZN(_032_)
);

NAND2_X1 _216_ (
  .A1(_059_),
  .A2(_032_),
  .ZN(_033_)
);

NAND2_X1 _217_ (
  .A1(_033_),
  .A2(_062_),
  .ZN(_034_)
);

AOI21_X1 _218_ (
  .A(_029_),
  .B1(_031_),
  .B2(_034_),
  .ZN(_008_)
);

AOI21_X1 _219_ (
  .A(_062_),
  .B1(_046_),
  .B2(_068_),
  .ZN(_035_)
);

NAND2_X1 _220_ (
  .A1(_023_),
  .A2(_035_),
  .ZN(_036_)
);

NOR2_X1 _221_ (
  .A1(_101_),
  .A2(_061_),
  .ZN(_037_)
);

NAND2_X1 _222_ (
  .A1(_025_),
  .A2(_037_),
  .ZN(_038_)
);

NAND3_X1 _223_ (
  .A1(_036_),
  .A2(_038_),
  .A3(_074_),
  .ZN(_039_)
);

NAND2_X1 _224_ (
  .A1(_076_),
  .A2(\coef[30] ),
  .ZN(_040_)
);

NAND2_X1 _225_ (
  .A1(_039_),
  .A2(_040_),
  .ZN(_009_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_117_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_116_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_115_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_114_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_113_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_112_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_111_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_110_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_109_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_108_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$a8d3b7b4edaf7d596a54a187c8ed4a9561fa625a\dctu

module \$paramod$adcdc49d3fc5249816d353bb65629f56cf0927d3\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X2 _069_ (
  .A(x[1]),
  .ZN(_008_)
);

NAND2_X4 _070_ (
  .A1(_008_),
  .A2(x[0]),
  .ZN(_009_)
);

INV_X2 _071_ (
  .A(x[0]),
  .ZN(_010_)
);

NAND2_X4 _072_ (
  .A1(_010_),
  .A2(x[1]),
  .ZN(_011_)
);

NAND2_X4 _073_ (
  .A1(_009_),
  .A2(_011_),
  .ZN(_012_)
);

INV_X1 _074_ (
  .A(y[0]),
  .ZN(_013_)
);

NAND2_X4 _075_ (
  .A1(_012_),
  .A2(_013_),
  .ZN(_014_)
);

NAND3_X4 _076_ (
  .A1(_009_),
  .A2(_011_),
  .A3(y[0]),
  .ZN(_015_)
);

NAND2_X4 _077_ (
  .A1(_014_),
  .A2(_015_),
  .ZN(_016_)
);

BUF_X4 _078_ (
  .A(y[1]),
  .Z(_017_)
);

INV_X2 _079_ (
  .A(_017_),
  .ZN(_018_)
);

NAND2_X4 _080_ (
  .A1(_016_),
  .A2(_018_),
  .ZN(_019_)
);

NAND3_X2 _081_ (
  .A1(_014_),
  .A2(_015_),
  .A3(_017_),
  .ZN(_020_)
);

BUF_X1 _082_ (
  .A(y[2]),
  .Z(_021_)
);

NAND3_X1 _083_ (
  .A1(_019_),
  .A2(_020_),
  .A3(_021_),
  .ZN(_022_)
);

NAND3_X2 _084_ (
  .A1(_014_),
  .A2(_015_),
  .A3(_018_),
  .ZN(_023_)
);

NAND3_X1 _085_ (
  .A1(_009_),
  .A2(_011_),
  .A3(_013_),
  .ZN(_024_)
);

NAND2_X1 _086_ (
  .A1(_008_),
  .A2(_010_),
  .ZN(_025_)
);

NAND2_X1 _087_ (
  .A1(x[1]),
  .A2(x[0]),
  .ZN(_026_)
);

NAND3_X1 _088_ (
  .A1(_025_),
  .A2(y[0]),
  .A3(_026_),
  .ZN(_027_)
);

NAND3_X1 _089_ (
  .A1(_024_),
  .A2(_027_),
  .A3(_017_),
  .ZN(_028_)
);

INV_X1 _090_ (
  .A(_021_),
  .ZN(_029_)
);

NAND3_X1 _091_ (
  .A1(_023_),
  .A2(_028_),
  .A3(_029_),
  .ZN(_030_)
);

CLKBUF_X3 _092_ (
  .A(ena),
  .Z(_031_)
);

NAND3_X1 _093_ (
  .A1(_022_),
  .A2(_030_),
  .A3(_031_),
  .ZN(_032_)
);

INV_X1 _094_ (
  .A(_031_),
  .ZN(_033_)
);

NAND2_X1 _095_ (
  .A1(_033_),
  .A2(\coef[21] ),
  .ZN(_034_)
);

NAND2_X1 _096_ (
  .A1(_032_),
  .A2(_034_),
  .ZN(_000_)
);

NAND2_X1 _097_ (
  .A1(_012_),
  .A2(_018_),
  .ZN(_035_)
);

NAND3_X2 _098_ (
  .A1(_020_),
  .A2(_029_),
  .A3(_035_),
  .ZN(_036_)
);

INV_X2 _099_ (
  .A(_012_),
  .ZN(_037_)
);

NAND2_X4 _100_ (
  .A1(_037_),
  .A2(_017_),
  .ZN(_038_)
);

NAND3_X2 _101_ (
  .A1(_023_),
  .A2(_021_),
  .A3(_038_),
  .ZN(_039_)
);

NAND3_X1 _102_ (
  .A1(_036_),
  .A2(_039_),
  .A3(_031_),
  .ZN(_040_)
);

NAND2_X1 _103_ (
  .A1(_033_),
  .A2(\coef[22] ),
  .ZN(_041_)
);

NAND2_X1 _104_ (
  .A1(_040_),
  .A2(_041_),
  .ZN(_001_)
);

NAND3_X1 _105_ (
  .A1(_019_),
  .A2(_029_),
  .A3(_038_),
  .ZN(_042_)
);

NAND3_X1 _106_ (
  .A1(_028_),
  .A2(_021_),
  .A3(_035_),
  .ZN(_043_)
);

NAND3_X1 _107_ (
  .A1(_042_),
  .A2(_043_),
  .A3(_031_),
  .ZN(_044_)
);

NAND2_X1 _108_ (
  .A1(_033_),
  .A2(\coef[23] ),
  .ZN(_045_)
);

NAND2_X1 _109_ (
  .A1(_044_),
  .A2(_045_),
  .ZN(_002_)
);

NAND2_X2 _110_ (
  .A1(_036_),
  .A2(_039_),
  .ZN(_046_)
);

NAND2_X2 _111_ (
  .A1(_046_),
  .A2(_031_),
  .ZN(_047_)
);

NAND2_X1 _112_ (
  .A1(_033_),
  .A2(\coef[14] ),
  .ZN(_048_)
);

NAND2_X2 _113_ (
  .A1(_047_),
  .A2(_048_),
  .ZN(_003_)
);

NOR2_X1 _114_ (
  .A1(_031_),
  .A2(\coef[13] ),
  .ZN(_049_)
);

AOI21_X1 _115_ (
  .A(_049_),
  .B1(_016_),
  .B2(_031_),
  .ZN(_004_)
);

NAND2_X1 _116_ (
  .A1(_037_),
  .A2(_018_),
  .ZN(_050_)
);

NAND2_X1 _117_ (
  .A1(_012_),
  .A2(_017_),
  .ZN(_051_)
);

NAND2_X1 _118_ (
  .A1(_050_),
  .A2(_051_),
  .ZN(_052_)
);

MUX2_X2 _119_ (
  .A(\coef[28] ),
  .B(_052_),
  .S(_031_),
  .Z(_005_)
);

NAND3_X1 _120_ (
  .A1(_019_),
  .A2(_021_),
  .A3(_038_),
  .ZN(_053_)
);

NAND3_X1 _121_ (
  .A1(_028_),
  .A2(_029_),
  .A3(_035_),
  .ZN(_054_)
);

NAND3_X1 _122_ (
  .A1(_053_),
  .A2(_054_),
  .A3(_031_),
  .ZN(_055_)
);

NAND2_X1 _123_ (
  .A1(_033_),
  .A2(\coef[15] ),
  .ZN(_056_)
);

NAND2_X1 _124_ (
  .A1(_055_),
  .A2(_056_),
  .ZN(_006_)
);

NAND3_X1 _125_ (
  .A1(_019_),
  .A2(_029_),
  .A3(_051_),
  .ZN(_057_)
);

NAND3_X1 _126_ (
  .A1(_028_),
  .A2(_021_),
  .A3(_050_),
  .ZN(_058_)
);

NAND3_X1 _127_ (
  .A1(_057_),
  .A2(_058_),
  .A3(_031_),
  .ZN(_059_)
);

NAND2_X1 _128_ (
  .A1(_033_),
  .A2(\coef[12] ),
  .ZN(_060_)
);

NAND2_X1 _129_ (
  .A1(_059_),
  .A2(_060_),
  .ZN(_007_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_068_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_067_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_066_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_065_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_064_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_063_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_062_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_061_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$adcdc49d3fc5249816d353bb65629f56cf0927d3\dctu

module \$paramod$b266e2f77428397c53d4afd55bef1da32efe03d9\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _092_ (
  .A(x[0]),
  .ZN(_074_)
);

INV_X1 _093_ (
  .A(x[1]),
  .ZN(_075_)
);

BUF_X4 _094_ (
  .A(y[0]),
  .Z(_009_)
);

BUF_X4 _095_ (
  .A(y[1]),
  .Z(_010_)
);

XNOR2_X2 _096_ (
  .A(_009_),
  .B(_010_),
  .ZN(_011_)
);

INV_X1 _097_ (
  .A(_011_),
  .ZN(_012_)
);

BUF_X4 _098_ (
  .A(x[2]),
  .Z(_013_)
);

INV_X2 _099_ (
  .A(_013_),
  .ZN(_014_)
);

NAND2_X1 _100_ (
  .A1(_014_),
  .A2(_090_),
  .ZN(_015_)
);

OR2_X1 _101_ (
  .A1(_014_),
  .A2(_076_),
  .ZN(_016_)
);

NAND3_X1 _102_ (
  .A1(_012_),
  .A2(_015_),
  .A3(_016_),
  .ZN(_017_)
);

OR2_X1 _103_ (
  .A1(_088_),
  .A2(_013_),
  .ZN(_018_)
);

NAND2_X1 _104_ (
  .A1(_078_),
  .A2(_013_),
  .ZN(_019_)
);

NAND3_X1 _105_ (
  .A1(_011_),
  .A2(_018_),
  .A3(_019_),
  .ZN(_020_)
);

BUF_X1 _106_ (
  .A(ena),
  .Z(_021_)
);

NAND3_X1 _107_ (
  .A1(_017_),
  .A2(_020_),
  .A3(_021_),
  .ZN(_022_)
);

INV_X1 _108_ (
  .A(ena),
  .ZN(_023_)
);

NAND2_X1 _109_ (
  .A1(_023_),
  .A2(\coef[21] ),
  .ZN(_024_)
);

NAND2_X1 _110_ (
  .A1(_022_),
  .A2(_024_),
  .ZN(_000_)
);

NAND2_X1 _111_ (
  .A1(_014_),
  .A2(_077_),
  .ZN(_025_)
);

INV_X1 _112_ (
  .A(_077_),
  .ZN(_026_)
);

NAND2_X1 _113_ (
  .A1(_026_),
  .A2(_013_),
  .ZN(_027_)
);

INV_X1 _114_ (
  .A(_009_),
  .ZN(_028_)
);

NAND3_X1 _115_ (
  .A1(_025_),
  .A2(_027_),
  .A3(_028_),
  .ZN(_029_)
);

NAND2_X1 _116_ (
  .A1(_014_),
  .A2(_026_),
  .ZN(_030_)
);

NAND2_X1 _117_ (
  .A1(_013_),
  .A2(_077_),
  .ZN(_031_)
);

NAND3_X1 _118_ (
  .A1(_030_),
  .A2(_009_),
  .A3(_031_),
  .ZN(_032_)
);

INV_X1 _119_ (
  .A(_010_),
  .ZN(_033_)
);

NAND3_X1 _120_ (
  .A1(_029_),
  .A2(_032_),
  .A3(_033_),
  .ZN(_034_)
);

NAND3_X1 _121_ (
  .A1(_025_),
  .A2(_027_),
  .A3(_009_),
  .ZN(_035_)
);

NAND3_X1 _122_ (
  .A1(_030_),
  .A2(_028_),
  .A3(_031_),
  .ZN(_036_)
);

NAND3_X1 _123_ (
  .A1(_035_),
  .A2(_036_),
  .A3(_010_),
  .ZN(_037_)
);

NAND3_X1 _124_ (
  .A1(_034_),
  .A2(_037_),
  .A3(_021_),
  .ZN(_038_)
);

NAND2_X1 _125_ (
  .A1(_023_),
  .A2(\coef[22] ),
  .ZN(_039_)
);

NAND2_X1 _126_ (
  .A1(_038_),
  .A2(_039_),
  .ZN(_001_)
);

NOR2_X1 _127_ (
  .A1(_021_),
  .A2(\coef[23] ),
  .ZN(_040_)
);

XNOR2_X1 _128_ (
  .A(_011_),
  .B(_074_),
  .ZN(_041_)
);

AOI21_X2 _129_ (
  .A(_040_),
  .B1(_041_),
  .B2(_021_),
  .ZN(_002_)
);

NAND3_X1 _130_ (
  .A1(_035_),
  .A2(_036_),
  .A3(_033_),
  .ZN(_042_)
);

NAND3_X1 _131_ (
  .A1(_029_),
  .A2(_032_),
  .A3(_010_),
  .ZN(_043_)
);

NAND3_X1 _132_ (
  .A1(_042_),
  .A2(_043_),
  .A3(_021_),
  .ZN(_044_)
);

NAND2_X1 _133_ (
  .A1(_023_),
  .A2(\coef[14] ),
  .ZN(_045_)
);

NAND2_X1 _134_ (
  .A1(_044_),
  .A2(_045_),
  .ZN(_003_)
);

NAND2_X1 _135_ (
  .A1(_014_),
  .A2(_086_),
  .ZN(_046_)
);

OR2_X1 _136_ (
  .A1(_014_),
  .A2(_080_),
  .ZN(_047_)
);

NAND3_X1 _137_ (
  .A1(_012_),
  .A2(_046_),
  .A3(_047_),
  .ZN(_048_)
);

INV_X1 _138_ (
  .A(_084_),
  .ZN(_049_)
);

NAND2_X1 _139_ (
  .A1(_014_),
  .A2(_049_),
  .ZN(_050_)
);

NAND2_X1 _140_ (
  .A1(_013_),
  .A2(_082_),
  .ZN(_051_)
);

NAND3_X1 _141_ (
  .A1(_011_),
  .A2(_050_),
  .A3(_051_),
  .ZN(_052_)
);

NAND3_X1 _142_ (
  .A1(_048_),
  .A2(_052_),
  .A3(_021_),
  .ZN(_053_)
);

NAND2_X1 _143_ (
  .A1(_023_),
  .A2(\coef[13] ),
  .ZN(_054_)
);

NAND2_X1 _144_ (
  .A1(_053_),
  .A2(_054_),
  .ZN(_004_)
);

NOR2_X1 _145_ (
  .A1(_013_),
  .A2(_080_),
  .ZN(_055_)
);

AOI21_X1 _146_ (
  .A(_055_),
  .B1(_086_),
  .B2(_013_),
  .ZN(_056_)
);

NAND2_X1 _147_ (
  .A1(_056_),
  .A2(_012_),
  .ZN(_057_)
);

NAND2_X1 _148_ (
  .A1(_049_),
  .A2(_013_),
  .ZN(_058_)
);

NAND2_X1 _149_ (
  .A1(_014_),
  .A2(_082_),
  .ZN(_059_)
);

NAND3_X1 _150_ (
  .A1(_011_),
  .A2(_058_),
  .A3(_059_),
  .ZN(_060_)
);

NAND3_X1 _151_ (
  .A1(_057_),
  .A2(_021_),
  .A3(_060_),
  .ZN(_061_)
);

NAND2_X1 _152_ (
  .A1(_023_),
  .A2(\coef[28] ),
  .ZN(_062_)
);

NAND2_X1 _153_ (
  .A1(_061_),
  .A2(_062_),
  .ZN(_005_)
);

NOR2_X1 _154_ (
  .A1(_021_),
  .A2(\coef[15] ),
  .ZN(_063_)
);

XNOR2_X1 _155_ (
  .A(_011_),
  .B(x[1]),
  .ZN(_064_)
);

AOI21_X2 _156_ (
  .A(_063_),
  .B1(_064_),
  .B2(_021_),
  .ZN(_006_)
);

NOR2_X1 _157_ (
  .A1(ena),
  .A2(\coef[12] ),
  .ZN(_065_)
);

XNOR2_X1 _158_ (
  .A(_011_),
  .B(_014_),
  .ZN(_008_)
);

AOI21_X2 _159_ (
  .A(_065_),
  .B1(_008_),
  .B2(_021_),
  .ZN(_007_)
);

HA_X1 _160_ (
  .A(_074_),
  .B(_075_),
  .CO(_076_),
  .S(_077_)
);

HA_X1 _161_ (
  .A(_074_),
  .B(_075_),
  .CO(_078_),
  .S(_079_)
);

HA_X1 _162_ (
  .A(_074_),
  .B(x[1]),
  .CO(_080_),
  .S(_081_)
);

HA_X1 _163_ (
  .A(_074_),
  .B(x[1]),
  .CO(_082_),
  .S(_083_)
);

HA_X1 _164_ (
  .A(x[0]),
  .B(_075_),
  .CO(_084_),
  .S(_085_)
);

HA_X1 _165_ (
  .A(x[0]),
  .B(_075_),
  .CO(_086_),
  .S(_087_)
);

HA_X1 _166_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_088_),
  .S(_089_)
);

HA_X1 _167_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_090_),
  .S(_091_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_073_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_072_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_071_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_070_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_069_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_068_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_067_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_066_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$b266e2f77428397c53d4afd55bef1da32efe03d9\dctu

module \$paramod$b53123087aafc52fe604e5dcf6b6b1b8d73b2231\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _054_ (
  .A(x[1]),
  .ZN(_004_)
);

INV_X2 _055_ (
  .A(x[2]),
  .ZN(_005_)
);

NAND2_X2 _056_ (
  .A1(_004_),
  .A2(_005_),
  .ZN(_006_)
);

INV_X1 _057_ (
  .A(y[0]),
  .ZN(_007_)
);

NAND2_X1 _058_ (
  .A1(x[1]),
  .A2(x[2]),
  .ZN(_008_)
);

NAND3_X1 _059_ (
  .A1(_006_),
  .A2(_007_),
  .A3(_008_),
  .ZN(_009_)
);

INV_X1 _060_ (
  .A(x[0]),
  .ZN(_010_)
);

NAND2_X2 _061_ (
  .A1(_005_),
  .A2(_010_),
  .ZN(_011_)
);

NAND2_X1 _062_ (
  .A1(x[2]),
  .A2(x[0]),
  .ZN(_012_)
);

NAND3_X2 _063_ (
  .A1(_011_),
  .A2(y[0]),
  .A3(_012_),
  .ZN(_013_)
);

NAND2_X1 _064_ (
  .A1(_009_),
  .A2(_013_),
  .ZN(_014_)
);

CLKBUF_X2 _065_ (
  .A(y[1]),
  .Z(_015_)
);

INV_X1 _066_ (
  .A(_015_),
  .ZN(_016_)
);

NAND2_X1 _067_ (
  .A1(_014_),
  .A2(_016_),
  .ZN(_017_)
);

NAND3_X1 _068_ (
  .A1(_011_),
  .A2(_007_),
  .A3(_012_),
  .ZN(_018_)
);

NAND3_X2 _069_ (
  .A1(_006_),
  .A2(y[0]),
  .A3(_008_),
  .ZN(_019_)
);

NAND3_X1 _070_ (
  .A1(_018_),
  .A2(_019_),
  .A3(_015_),
  .ZN(_020_)
);

CLKBUF_X2 _071_ (
  .A(y[2]),
  .Z(_021_)
);

INV_X1 _072_ (
  .A(_021_),
  .ZN(_022_)
);

NAND3_X1 _073_ (
  .A1(_017_),
  .A2(_020_),
  .A3(_022_),
  .ZN(_023_)
);

NAND2_X1 _074_ (
  .A1(_018_),
  .A2(_019_),
  .ZN(_024_)
);

NAND2_X1 _075_ (
  .A1(_024_),
  .A2(_015_),
  .ZN(_025_)
);

NAND3_X1 _076_ (
  .A1(_009_),
  .A2(_013_),
  .A3(_016_),
  .ZN(_026_)
);

NAND3_X1 _077_ (
  .A1(_025_),
  .A2(_026_),
  .A3(_021_),
  .ZN(_027_)
);

BUF_X2 _078_ (
  .A(ena),
  .Z(_028_)
);

NAND3_X1 _079_ (
  .A1(_023_),
  .A2(_027_),
  .A3(_028_),
  .ZN(_029_)
);

INV_X1 _080_ (
  .A(_028_),
  .ZN(_030_)
);

NAND2_X1 _081_ (
  .A1(_030_),
  .A2(\coef[13] ),
  .ZN(_031_)
);

NAND2_X1 _082_ (
  .A1(_029_),
  .A2(_031_),
  .ZN(_000_)
);

NAND3_X1 _083_ (
  .A1(_017_),
  .A2(_020_),
  .A3(_021_),
  .ZN(_032_)
);

NAND3_X1 _084_ (
  .A1(_025_),
  .A2(_026_),
  .A3(_022_),
  .ZN(_033_)
);

NAND3_X1 _085_ (
  .A1(_032_),
  .A2(_033_),
  .A3(_028_),
  .ZN(_034_)
);

NAND2_X1 _086_ (
  .A1(_030_),
  .A2(\coef[10] ),
  .ZN(_035_)
);

NAND2_X1 _087_ (
  .A1(_034_),
  .A2(_035_),
  .ZN(_001_)
);

NAND2_X1 _088_ (
  .A1(_011_),
  .A2(_012_),
  .ZN(_036_)
);

NAND2_X1 _089_ (
  .A1(_036_),
  .A2(_007_),
  .ZN(_037_)
);

NAND3_X1 _090_ (
  .A1(_037_),
  .A2(_019_),
  .A3(_016_),
  .ZN(_038_)
);

NAND2_X2 _091_ (
  .A1(_006_),
  .A2(_008_),
  .ZN(_039_)
);

NAND2_X2 _092_ (
  .A1(_039_),
  .A2(_007_),
  .ZN(_040_)
);

NAND3_X2 _093_ (
  .A1(_040_),
  .A2(_013_),
  .A3(_015_),
  .ZN(_041_)
);

NAND2_X1 _094_ (
  .A1(_038_),
  .A2(_041_),
  .ZN(_042_)
);

NAND2_X1 _095_ (
  .A1(_042_),
  .A2(_022_),
  .ZN(_043_)
);

NAND3_X1 _096_ (
  .A1(_038_),
  .A2(_041_),
  .A3(_021_),
  .ZN(_044_)
);

NAND3_X1 _097_ (
  .A1(_043_),
  .A2(_044_),
  .A3(_028_),
  .ZN(_045_)
);

NAND2_X1 _098_ (
  .A1(_030_),
  .A2(\coef[29] ),
  .ZN(_046_)
);

NAND2_X1 _099_ (
  .A1(_045_),
  .A2(_046_),
  .ZN(_002_)
);

NOR2_X1 _100_ (
  .A1(_028_),
  .A2(\coef[30] ),
  .ZN(_047_)
);

XNOR2_X1 _101_ (
  .A(_015_),
  .B(_021_),
  .ZN(_048_)
);

XNOR2_X1 _102_ (
  .A(_048_),
  .B(_039_),
  .ZN(_049_)
);

AOI21_X1 _103_ (
  .A(_047_),
  .B1(_049_),
  .B2(_028_),
  .ZN(_003_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_053_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_052_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_051_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_050_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[10] , \coef[13] , \coef[10] , \coef[10] , \coef[13] , \coef[10] , \coef[13] , \coef[10] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$b53123087aafc52fe604e5dcf6b6b1b8d73b2231\dctu

module \$paramod$141303f1e6ff0436e3fa44dd8e1d8f51afed9a78\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _069_ (
  .A(y[0]),
  .ZN(_051_)
);

INV_X1 _070_ (
  .A(y[1]),
  .ZN(_052_)
);

BUF_X4 _071_ (
  .A(ena),
  .Z(_008_)
);

INV_X4 _072_ (
  .A(_008_),
  .ZN(_009_)
);

NAND2_X1 _073_ (
  .A1(_009_),
  .A2(\coef[13] ),
  .ZN(_010_)
);

BUF_X4 _074_ (
  .A(y[2]),
  .Z(_011_)
);

INV_X4 _075_ (
  .A(_011_),
  .ZN(_012_)
);

OAI21_X1 _076_ (
  .A(_010_),
  .B1(_012_),
  .B2(_009_),
  .ZN(_000_)
);

INV_X1 _077_ (
  .A(_055_),
  .ZN(_013_)
);

NAND2_X1 _078_ (
  .A1(_013_),
  .A2(_011_),
  .ZN(_014_)
);

NAND2_X1 _079_ (
  .A1(_012_),
  .A2(_065_),
  .ZN(_015_)
);

NAND3_X1 _080_ (
  .A1(_014_),
  .A2(_015_),
  .A3(_008_),
  .ZN(_016_)
);

NAND2_X1 _081_ (
  .A1(_009_),
  .A2(\coef[14] ),
  .ZN(_017_)
);

NAND2_X1 _082_ (
  .A1(_016_),
  .A2(_017_),
  .ZN(_001_)
);

INV_X1 _083_ (
  .A(_063_),
  .ZN(_018_)
);

NAND2_X1 _084_ (
  .A1(_018_),
  .A2(_011_),
  .ZN(_019_)
);

NAND2_X1 _085_ (
  .A1(_012_),
  .A2(_057_),
  .ZN(_020_)
);

NAND3_X1 _086_ (
  .A1(_019_),
  .A2(_020_),
  .A3(_008_),
  .ZN(_021_)
);

NAND2_X1 _087_ (
  .A1(_009_),
  .A2(\coef[15] ),
  .ZN(_022_)
);

NAND2_X1 _088_ (
  .A1(_021_),
  .A2(_022_),
  .ZN(_002_)
);

INV_X1 _089_ (
  .A(_067_),
  .ZN(_023_)
);

NAND2_X1 _090_ (
  .A1(_023_),
  .A2(_011_),
  .ZN(_024_)
);

NAND2_X1 _091_ (
  .A1(_012_),
  .A2(_053_),
  .ZN(_025_)
);

NAND3_X1 _092_ (
  .A1(_024_),
  .A2(_025_),
  .A3(_008_),
  .ZN(_026_)
);

NAND2_X1 _093_ (
  .A1(_009_),
  .A2(\coef[12] ),
  .ZN(_027_)
);

NAND2_X1 _094_ (
  .A1(_026_),
  .A2(_027_),
  .ZN(_003_)
);

NAND2_X1 _095_ (
  .A1(_009_),
  .A2(\coef[21] ),
  .ZN(_028_)
);

OAI21_X1 _096_ (
  .A(_028_),
  .B1(y[1]),
  .B2(_009_),
  .ZN(_004_)
);

NAND2_X1 _097_ (
  .A1(_009_),
  .A2(\coef[22] ),
  .ZN(_029_)
);

NAND2_X1 _098_ (
  .A1(_011_),
  .A2(_053_),
  .ZN(_030_)
);

NAND2_X1 _099_ (
  .A1(_030_),
  .A2(_008_),
  .ZN(_031_)
);

NOR2_X1 _100_ (
  .A1(_067_),
  .A2(_011_),
  .ZN(_032_)
);

OAI21_X1 _101_ (
  .A(_029_),
  .B1(_031_),
  .B2(_032_),
  .ZN(_005_)
);

INV_X1 _102_ (
  .A(_059_),
  .ZN(_033_)
);

NAND2_X1 _103_ (
  .A1(_033_),
  .A2(_011_),
  .ZN(_034_)
);

NAND2_X1 _104_ (
  .A1(_012_),
  .A2(_061_),
  .ZN(_035_)
);

NAND3_X1 _105_ (
  .A1(_034_),
  .A2(_035_),
  .A3(_008_),
  .ZN(_036_)
);

NAND2_X1 _106_ (
  .A1(_009_),
  .A2(\coef[23] ),
  .ZN(_037_)
);

NAND2_X1 _107_ (
  .A1(_036_),
  .A2(_037_),
  .ZN(_006_)
);

INV_X1 _108_ (
  .A(_054_),
  .ZN(_038_)
);

NAND2_X1 _109_ (
  .A1(_012_),
  .A2(_038_),
  .ZN(_039_)
);

NAND2_X1 _110_ (
  .A1(_011_),
  .A2(_054_),
  .ZN(_040_)
);

NAND3_X1 _111_ (
  .A1(_039_),
  .A2(_008_),
  .A3(_040_),
  .ZN(_041_)
);

NAND2_X1 _112_ (
  .A1(_009_),
  .A2(\coef[28] ),
  .ZN(_042_)
);

NAND2_X1 _113_ (
  .A1(_041_),
  .A2(_042_),
  .ZN(_007_)
);

HA_X1 _114_ (
  .A(_051_),
  .B(_052_),
  .CO(_053_),
  .S(_054_)
);

HA_X1 _115_ (
  .A(_051_),
  .B(_052_),
  .CO(_055_),
  .S(_056_)
);

HA_X1 _116_ (
  .A(_051_),
  .B(y[1]),
  .CO(_057_),
  .S(_058_)
);

HA_X1 _117_ (
  .A(_051_),
  .B(y[1]),
  .CO(_059_),
  .S(_060_)
);

HA_X1 _118_ (
  .A(y[0]),
  .B(_052_),
  .CO(_061_),
  .S(_062_)
);

HA_X1 _119_ (
  .A(y[0]),
  .B(_052_),
  .CO(_063_),
  .S(_064_)
);

HA_X1 _120_ (
  .A(y[0]),
  .B(y[1]),
  .CO(_065_),
  .S(_066_)
);

HA_X1 _121_ (
  .A(y[0]),
  .B(y[1]),
  .CO(_067_),
  .S(_068_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_046_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_045_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_044_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_049_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_050_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_043_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_048_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_047_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$141303f1e6ff0436e3fa44dd8e1d8f51afed9a78\dctu

module jpeg_rle(input clk, input rst, input ena, input dstrb, input [11:0] din, output [3:0] size,
 output [3:0] rlen, output [11:0] amp, output douten, output bstart);
wire _0_;
wire ddstrb;
wire \rle_amp[0] ;
wire \rle_amp[10] ;
wire \rle_amp[11] ;
wire \rle_amp[1] ;
wire \rle_amp[2] ;
wire \rle_amp[3] ;
wire \rle_amp[4] ;
wire \rle_amp[5] ;
wire \rle_amp[6] ;
wire \rle_amp[7] ;
wire \rle_amp[8] ;
wire \rle_amp[9] ;
wire rle_dc;
wire rle_den;
wire \rle_rlen[0] ;
wire \rle_rlen[1] ;
wire \rle_rlen[2] ;
wire \rle_rlen[3] ;
wire \rle_size[0] ;
wire \rle_size[1] ;
wire \rle_size[2] ;
wire \rle_size[3] ;
wire \rz1_amp[0] ;
wire \rz1_amp[10] ;
wire \rz1_amp[11] ;
wire \rz1_amp[1] ;
wire \rz1_amp[2] ;
wire \rz1_amp[3] ;
wire \rz1_amp[4] ;
wire \rz1_amp[5] ;
wire \rz1_amp[6] ;
wire \rz1_amp[7] ;
wire \rz1_amp[8] ;
wire \rz1_amp[9] ;
wire rz1_dc;
wire rz1_den;
wire \rz1_rlen[0] ;
wire \rz1_rlen[1] ;
wire \rz1_rlen[2] ;
wire \rz1_rlen[3] ;
wire \rz1_size[0] ;
wire \rz1_size[1] ;
wire \rz1_size[2] ;
wire \rz1_size[3] ;
wire \rz2_amp[0] ;
wire \rz2_amp[10] ;
wire \rz2_amp[11] ;
wire \rz2_amp[1] ;
wire \rz2_amp[2] ;
wire \rz2_amp[3] ;
wire \rz2_amp[4] ;
wire \rz2_amp[5] ;
wire \rz2_amp[6] ;
wire \rz2_amp[7] ;
wire \rz2_amp[8] ;
wire \rz2_amp[9] ;
wire rz2_dc;
wire rz2_den;
wire \rz2_rlen[0] ;
wire \rz2_rlen[1] ;
wire \rz2_rlen[2] ;
wire \rz2_rlen[3] ;
wire \rz2_size[0] ;
wire \rz2_size[1] ;
wire \rz2_size[2] ;
wire \rz2_size[3] ;
wire \rz3_amp[0] ;
wire \rz3_amp[10] ;
wire \rz3_amp[11] ;
wire \rz3_amp[1] ;
wire \rz3_amp[2] ;
wire \rz3_amp[3] ;
wire \rz3_amp[4] ;
wire \rz3_amp[5] ;
wire \rz3_amp[6] ;
wire \rz3_amp[7] ;
wire \rz3_amp[8] ;
wire \rz3_amp[9] ;
wire rz3_dc;
wire rz3_den;
wire \rz3_rlen[0] ;
wire \rz3_rlen[1] ;
wire \rz3_rlen[2] ;
wire \rz3_rlen[3] ;
wire \rz3_size[0] ;
wire \rz3_size[1] ;
wire \rz3_size[2] ;
wire \rz3_size[3] ;

DFF_X1 ddstrb$_DFF_P_ (
  .D(dstrb),
  .CK(clk),
  .Q(ddstrb),
  .QN(_0_)
);

jpeg_rle1 rle (
  .clk(clk),
  .rst(rst),
  .ena(ena),
  .go(ddstrb),
  .din(din),
  .rlen({\rle_rlen[3] , \rle_rlen[2] , \rle_rlen[1] , \rle_rlen[0] }),
  .size({\rle_size[3] , \rle_size[2] , \rle_size[1] , \rle_size[0] }),
  .amp({\rle_amp[11] , \rle_amp[10] , \rle_amp[9] , \rle_amp[8] , \rle_amp[7] , \rle_amp[6] , \rle_amp[5] , \rle_amp[4] , \rle_amp[3] , \rle_amp[2] , \rle_amp[1] , \rle_amp[0] }),
  .den(rle_den),
  .dcterm(rle_dc)
);

jpeg_rzs_clone_498 rz1 (
  .clk(clk),
  .ena(ena),
  .rst(rst),
  .deni(rle_den),
  .dci(rle_dc),
  .rleni({\rle_rlen[3] , \rle_rlen[2] , \rle_rlen[1] , \rle_rlen[0] }),
  .sizei({\rle_size[3] , \rle_size[2] , \rle_size[1] , \rle_size[0] }),
  .ampi({\rle_amp[11] , \rle_amp[10] , \rle_amp[9] , \rle_amp[8] , \rle_amp[7] , \rle_amp[6] , \rle_amp[5] , \rle_amp[4] , \rle_amp[3] , \rle_amp[2] , \rle_amp[1] , \rle_amp[0] }),
  .deno(rz1_den),
  .dco(rz1_dc),
  .rleno({\rz1_rlen[3] , \rz1_rlen[2] , \rz1_rlen[1] , \rz1_rlen[0] }),
  .sizeo({\rz1_size[3] , \rz1_size[2] , \rz1_size[1] , \rz1_size[0] }),
  .ampo({\rz1_amp[11] , \rz1_amp[10] , \rz1_amp[9] , \rz1_amp[8] , \rz1_amp[7] , \rz1_amp[6] , \rz1_amp[5] , \rz1_amp[4] , \rz1_amp[3] , \rz1_amp[2] , \rz1_amp[1] , \rz1_amp[0] })
);

jpeg_rzs rz2 (
  .clk(clk),
  .ena(ena),
  .rst(rst),
  .deni(rz1_den),
  .dci(rz1_dc),
  .rleni({\rz1_rlen[3] , \rz1_rlen[2] , \rz1_rlen[1] , \rz1_rlen[0] }),
  .sizei({\rz1_size[3] , \rz1_size[2] , \rz1_size[1] , \rz1_size[0] }),
  .ampi({\rz1_amp[11] , \rz1_amp[10] , \rz1_amp[9] , \rz1_amp[8] , \rz1_amp[7] , \rz1_amp[6] , \rz1_amp[5] , \rz1_amp[4] , \rz1_amp[3] , \rz1_amp[2] , \rz1_amp[1] , \rz1_amp[0] }),
  .deno(rz2_den),
  .dco(rz2_dc),
  .rleno({\rz2_rlen[3] , \rz2_rlen[2] , \rz2_rlen[1] , \rz2_rlen[0] }),
  .sizeo({\rz2_size[3] , \rz2_size[2] , \rz2_size[1] , \rz2_size[0] }),
  .ampo({\rz2_amp[11] , \rz2_amp[10] , \rz2_amp[9] , \rz2_amp[8] , \rz2_amp[7] , \rz2_amp[6] , \rz2_amp[5] , \rz2_amp[4] , \rz2_amp[3] , \rz2_amp[2] , \rz2_amp[1] , \rz2_amp[0] })
);

jpeg_rzs rz3 (
  .clk(clk),
  .ena(ena),
  .rst(rst),
  .deni(rz2_den),
  .dci(rz2_dc),
  .rleni({\rz2_rlen[3] , \rz2_rlen[2] , \rz2_rlen[1] , \rz2_rlen[0] }),
  .sizei({\rz2_size[3] , \rz2_size[2] , \rz2_size[1] , \rz2_size[0] }),
  .ampi({\rz2_amp[11] , \rz2_amp[10] , \rz2_amp[9] , \rz2_amp[8] , \rz2_amp[7] , \rz2_amp[6] , \rz2_amp[5] , \rz2_amp[4] , \rz2_amp[3] , \rz2_amp[2] , \rz2_amp[1] , \rz2_amp[0] }),
  .deno(rz3_den),
  .dco(rz3_dc),
  .rleno({\rz3_rlen[3] , \rz3_rlen[2] , \rz3_rlen[1] , \rz3_rlen[0] }),
  .sizeo({\rz3_size[3] , \rz3_size[2] , \rz3_size[1] , \rz3_size[0] }),
  .ampo({\rz3_amp[11] , \rz3_amp[10] , \rz3_amp[9] , \rz3_amp[8] , \rz3_amp[7] , \rz3_amp[6] , \rz3_amp[5] , \rz3_amp[4] , \rz3_amp[3] , \rz3_amp[2] , \rz3_amp[1] , \rz3_amp[0] })
);

jpeg_rzs_clone_94 rz4 (
  .clk(clk),
  .ena(ena),
  .rst(rst),
  .deni(rz3_den),
  .dci(rz3_dc),
  .rleni({\rz3_rlen[3] , \rz3_rlen[2] , \rz3_rlen[1] , \rz3_rlen[0] }),
  .sizei({\rz3_size[3] , \rz3_size[2] , \rz3_size[1] , \rz3_size[0] }),
  .ampi({\rz3_amp[11] , \rz3_amp[10] , \rz3_amp[9] , \rz3_amp[8] , \rz3_amp[7] , \rz3_amp[6] , \rz3_amp[5] , \rz3_amp[4] , \rz3_amp[3] , \rz3_amp[2] , \rz3_amp[1] , \rz3_amp[0] }),
  .deno(douten),
  .dco(bstart),
  .rleno(rlen),
  .sizeo(size),
  .ampo(amp)
);
endmodule //jpeg_rle

module \$paramod$bb43d9c07810ea45f23a5f680ee116bafcd9334e\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _063_ (
  .A(x[0]),
  .ZN(_049_)
);

INV_X1 _064_ (
  .A(x[1]),
  .ZN(_050_)
);

INV_X1 _065_ (
  .A(_052_),
  .ZN(_008_)
);

BUF_X4 _066_ (
  .A(x[2]),
  .Z(_009_)
);

NAND2_X1 _067_ (
  .A1(_008_),
  .A2(_009_),
  .ZN(_010_)
);

INV_X4 _068_ (
  .A(_009_),
  .ZN(_011_)
);

NAND2_X2 _069_ (
  .A1(_011_),
  .A2(_052_),
  .ZN(_012_)
);

BUF_X4 _070_ (
  .A(ena),
  .Z(_013_)
);

NAND3_X1 _071_ (
  .A1(_010_),
  .A2(_012_),
  .A3(_013_),
  .ZN(_014_)
);

INV_X4 _072_ (
  .A(_013_),
  .ZN(_015_)
);

NAND2_X1 _073_ (
  .A1(_015_),
  .A2(\coef[21] ),
  .ZN(_016_)
);

NAND2_X1 _074_ (
  .A1(_014_),
  .A2(_016_),
  .ZN(_000_)
);

NAND2_X1 _075_ (
  .A1(_015_),
  .A2(\coef[22] ),
  .ZN(_017_)
);

NAND2_X1 _076_ (
  .A1(_009_),
  .A2(_057_),
  .ZN(_018_)
);

NAND2_X1 _077_ (
  .A1(_018_),
  .A2(_013_),
  .ZN(_019_)
);

NOR2_X1 _078_ (
  .A1(_009_),
  .A2(_055_),
  .ZN(_020_)
);

OAI21_X1 _079_ (
  .A(_017_),
  .B1(_019_),
  .B2(_020_),
  .ZN(_001_)
);

INV_X1 _080_ (
  .A(_061_),
  .ZN(_021_)
);

NAND2_X1 _081_ (
  .A1(_021_),
  .A2(_009_),
  .ZN(_022_)
);

NAND2_X2 _082_ (
  .A1(_011_),
  .A2(_051_),
  .ZN(_023_)
);

NAND3_X1 _083_ (
  .A1(_022_),
  .A2(_023_),
  .A3(_013_),
  .ZN(_024_)
);

NAND2_X1 _084_ (
  .A1(_015_),
  .A2(\coef[23] ),
  .ZN(_025_)
);

NAND2_X1 _085_ (
  .A1(_024_),
  .A2(_025_),
  .ZN(_002_)
);

INV_X1 _086_ (
  .A(_059_),
  .ZN(_026_)
);

NAND2_X1 _087_ (
  .A1(_026_),
  .A2(_009_),
  .ZN(_027_)
);

NAND2_X2 _088_ (
  .A1(_011_),
  .A2(_053_),
  .ZN(_028_)
);

NAND3_X1 _089_ (
  .A1(_027_),
  .A2(_028_),
  .A3(_013_),
  .ZN(_029_)
);

NAND2_X1 _090_ (
  .A1(_015_),
  .A2(\coef[14] ),
  .ZN(_030_)
);

NAND2_X1 _091_ (
  .A1(_029_),
  .A2(_030_),
  .ZN(_003_)
);

NAND2_X1 _092_ (
  .A1(_015_),
  .A2(\coef[13] ),
  .ZN(_031_)
);

OAI21_X1 _093_ (
  .A(_031_),
  .B1(x[0]),
  .B2(_015_),
  .ZN(_004_)
);

NAND2_X1 _094_ (
  .A1(_015_),
  .A2(\coef[28] ),
  .ZN(_032_)
);

OAI21_X1 _095_ (
  .A(_032_),
  .B1(x[1]),
  .B2(_015_),
  .ZN(_005_)
);

NAND2_X1 _096_ (
  .A1(_015_),
  .A2(\coef[15] ),
  .ZN(_033_)
);

NAND2_X1 _097_ (
  .A1(_009_),
  .A2(_051_),
  .ZN(_034_)
);

NAND2_X1 _098_ (
  .A1(_034_),
  .A2(_013_),
  .ZN(_035_)
);

NOR2_X1 _099_ (
  .A1(_009_),
  .A2(_061_),
  .ZN(_036_)
);

OAI21_X1 _100_ (
  .A(_033_),
  .B1(_035_),
  .B2(_036_),
  .ZN(_006_)
);

NAND2_X1 _101_ (
  .A1(_015_),
  .A2(\coef[12] ),
  .ZN(_037_)
);

NAND2_X1 _102_ (
  .A1(_009_),
  .A2(_053_),
  .ZN(_038_)
);

NAND2_X1 _103_ (
  .A1(_038_),
  .A2(_013_),
  .ZN(_039_)
);

NOR2_X1 _104_ (
  .A1(_009_),
  .A2(_059_),
  .ZN(_040_)
);

OAI21_X1 _105_ (
  .A(_037_),
  .B1(_039_),
  .B2(_040_),
  .ZN(_007_)
);

HA_X1 _106_ (
  .A(_049_),
  .B(_050_),
  .CO(_051_),
  .S(_052_)
);

HA_X1 _107_ (
  .A(_049_),
  .B(x[1]),
  .CO(_053_),
  .S(_054_)
);

HA_X1 _108_ (
  .A(_049_),
  .B(x[1]),
  .CO(_055_),
  .S(_056_)
);

HA_X1 _109_ (
  .A(x[0]),
  .B(_050_),
  .CO(_057_),
  .S(_058_)
);

HA_X1 _110_ (
  .A(x[0]),
  .B(_050_),
  .CO(_059_),
  .S(_060_)
);

HA_X1 _111_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_061_),
  .S(_062_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_048_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_047_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_046_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_045_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_044_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_043_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_042_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_041_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$bb43d9c07810ea45f23a5f680ee116bafcd9334e\dctu

module \$paramod$bd585d540938973e77d9fdfafe68a3c54bf55cb8\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X2 _053_ (
  .A(x[2]),
  .ZN(_004_)
);

INV_X1 _054_ (
  .A(x[0]),
  .ZN(_005_)
);

NAND2_X2 _055_ (
  .A1(_004_),
  .A2(_005_),
  .ZN(_006_)
);

INV_X1 _056_ (
  .A(y[0]),
  .ZN(_007_)
);

NAND2_X1 _057_ (
  .A1(x[2]),
  .A2(x[0]),
  .ZN(_008_)
);

NAND3_X1 _058_ (
  .A1(_006_),
  .A2(_007_),
  .A3(_008_),
  .ZN(_009_)
);

INV_X1 _059_ (
  .A(x[1]),
  .ZN(_010_)
);

NAND2_X2 _060_ (
  .A1(_010_),
  .A2(_004_),
  .ZN(_011_)
);

NAND2_X1 _061_ (
  .A1(x[1]),
  .A2(x[2]),
  .ZN(_012_)
);

NAND3_X1 _062_ (
  .A1(_011_),
  .A2(y[0]),
  .A3(_012_),
  .ZN(_013_)
);

NAND2_X1 _063_ (
  .A1(_009_),
  .A2(_013_),
  .ZN(_014_)
);

NAND2_X1 _064_ (
  .A1(_014_),
  .A2(y[1]),
  .ZN(_015_)
);

NAND3_X1 _065_ (
  .A1(_011_),
  .A2(_007_),
  .A3(_012_),
  .ZN(_016_)
);

NAND3_X1 _066_ (
  .A1(_006_),
  .A2(y[0]),
  .A3(_008_),
  .ZN(_017_)
);

INV_X1 _067_ (
  .A(y[1]),
  .ZN(_018_)
);

NAND3_X1 _068_ (
  .A1(_016_),
  .A2(_017_),
  .A3(_018_),
  .ZN(_019_)
);

BUF_X1 _069_ (
  .A(y[2]),
  .Z(_020_)
);

INV_X1 _070_ (
  .A(_020_),
  .ZN(_021_)
);

NAND3_X1 _071_ (
  .A1(_015_),
  .A2(_019_),
  .A3(_021_),
  .ZN(_022_)
);

NAND2_X1 _072_ (
  .A1(_006_),
  .A2(_008_),
  .ZN(_023_)
);

NAND2_X1 _073_ (
  .A1(_023_),
  .A2(y[0]),
  .ZN(_024_)
);

NAND2_X1 _074_ (
  .A1(_011_),
  .A2(_012_),
  .ZN(_025_)
);

NAND2_X1 _075_ (
  .A1(_025_),
  .A2(_007_),
  .ZN(_026_)
);

NAND3_X1 _076_ (
  .A1(_024_),
  .A2(_026_),
  .A3(_018_),
  .ZN(_027_)
);

NAND3_X1 _077_ (
  .A1(_009_),
  .A2(_013_),
  .A3(y[1]),
  .ZN(_028_)
);

NAND3_X1 _078_ (
  .A1(_027_),
  .A2(_028_),
  .A3(_020_),
  .ZN(_029_)
);

BUF_X2 _079_ (
  .A(ena),
  .Z(_030_)
);

NAND3_X1 _080_ (
  .A1(_022_),
  .A2(_029_),
  .A3(_030_),
  .ZN(_031_)
);

INV_X1 _081_ (
  .A(_030_),
  .ZN(_032_)
);

NAND2_X1 _082_ (
  .A1(_032_),
  .A2(\coef[13] ),
  .ZN(_033_)
);

NAND2_X1 _083_ (
  .A1(_031_),
  .A2(_033_),
  .ZN(_000_)
);

NAND3_X1 _084_ (
  .A1(_015_),
  .A2(_019_),
  .A3(_020_),
  .ZN(_034_)
);

NAND3_X1 _085_ (
  .A1(_027_),
  .A2(_028_),
  .A3(_021_),
  .ZN(_035_)
);

NAND3_X1 _086_ (
  .A1(_034_),
  .A2(_035_),
  .A3(_030_),
  .ZN(_036_)
);

NAND2_X1 _087_ (
  .A1(_032_),
  .A2(\coef[10] ),
  .ZN(_037_)
);

NAND2_X1 _088_ (
  .A1(_036_),
  .A2(_037_),
  .ZN(_001_)
);

NAND2_X1 _089_ (
  .A1(_023_),
  .A2(_007_),
  .ZN(_038_)
);

NAND3_X1 _090_ (
  .A1(_038_),
  .A2(_013_),
  .A3(_018_),
  .ZN(_039_)
);

NAND3_X1 _091_ (
  .A1(_026_),
  .A2(_017_),
  .A3(y[1]),
  .ZN(_040_)
);

NAND2_X1 _092_ (
  .A1(_039_),
  .A2(_040_),
  .ZN(_041_)
);

NAND2_X1 _093_ (
  .A1(_041_),
  .A2(_020_),
  .ZN(_042_)
);

NAND3_X1 _094_ (
  .A1(_039_),
  .A2(_040_),
  .A3(_021_),
  .ZN(_043_)
);

NAND3_X1 _095_ (
  .A1(_042_),
  .A2(_043_),
  .A3(_030_),
  .ZN(_044_)
);

NAND2_X1 _096_ (
  .A1(_032_),
  .A2(\coef[29] ),
  .ZN(_045_)
);

NAND2_X1 _097_ (
  .A1(_044_),
  .A2(_045_),
  .ZN(_002_)
);

NOR2_X1 _098_ (
  .A1(_030_),
  .A2(\coef[30] ),
  .ZN(_046_)
);

NAND2_X1 _099_ (
  .A1(_024_),
  .A2(_009_),
  .ZN(_047_)
);

XNOR2_X1 _100_ (
  .A(_047_),
  .B(_020_),
  .ZN(_048_)
);

AOI21_X2 _101_ (
  .A(_046_),
  .B1(_048_),
  .B2(_030_),
  .ZN(_003_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_052_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_051_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_050_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_049_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[10] , \coef[13] , \coef[10] , \coef[10] , \coef[13] , \coef[10] , \coef[13] , \coef[10] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$bd585d540938973e77d9fdfafe68a3c54bf55cb8\dctu

module \$paramod$bd5d8b7ea001bd9da1e8d07da4940a1f4c75e6b0\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _11_ (
  .A(x[1]),
  .ZN(_04_)
);

INV_X1 _12_ (
  .A(x[0]),
  .ZN(_05_)
);

NAND2_X1 _13_ (
  .A1(_04_),
  .A2(_05_),
  .ZN(_06_)
);

NAND2_X1 _14_ (
  .A1(x[1]),
  .A2(x[0]),
  .ZN(_07_)
);

NAND3_X1 _15_ (
  .A1(_06_),
  .A2(ena),
  .A3(_07_),
  .ZN(_01_)
);

INV_X1 _16_ (
  .A(ena),
  .ZN(_02_)
);

NAND2_X1 _17_ (
  .A1(_02_),
  .A2(\coef[30] ),
  .ZN(_03_)
);

NAND2_X1 _18_ (
  .A1(_01_),
  .A2(_03_),
  .ZN(_00_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_08_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac_clone_80644  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , _09_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_}),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$bd5d8b7ea001bd9da1e8d07da4940a1f4c75e6b0\dctu

module \$paramod$bfc28a02cfebf191b4a982c9147f38f65a3f3469\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _190_ (
  .A(x[0]),
  .ZN(_172_)
);

INV_X1 _191_ (
  .A(x[1]),
  .ZN(_173_)
);

INV_X2 _192_ (
  .A(x[2]),
  .ZN(_103_)
);

INV_X1 _193_ (
  .A(_175_),
  .ZN(_104_)
);

NAND2_X1 _194_ (
  .A1(_103_),
  .A2(_104_),
  .ZN(_105_)
);

BUF_X4 _195_ (
  .A(x[2]),
  .Z(_106_)
);

NAND2_X4 _196_ (
  .A1(_106_),
  .A2(_175_),
  .ZN(_107_)
);

NAND2_X1 _197_ (
  .A1(_105_),
  .A2(_107_),
  .ZN(_108_)
);

BUF_X4 _198_ (
  .A(y[0]),
  .Z(_109_)
);

BUF_X4 _199_ (
  .A(_109_),
  .Z(_110_)
);

NAND2_X1 _200_ (
  .A1(_108_),
  .A2(_110_),
  .ZN(_111_)
);

BUF_X8 _201_ (
  .A(_103_),
  .Z(_112_)
);

NAND2_X4 _202_ (
  .A1(_112_),
  .A2(_174_),
  .ZN(_113_)
);

INV_X1 _203_ (
  .A(_188_),
  .ZN(_114_)
);

NAND2_X1 _204_ (
  .A1(_114_),
  .A2(_106_),
  .ZN(_115_)
);

INV_X4 _205_ (
  .A(_109_),
  .ZN(_116_)
);

NAND3_X2 _206_ (
  .A1(_113_),
  .A2(_115_),
  .A3(_116_),
  .ZN(_117_)
);

NAND2_X1 _207_ (
  .A1(_111_),
  .A2(_117_),
  .ZN(_118_)
);

BUF_X4 _208_ (
  .A(y[1]),
  .Z(_119_)
);

BUF_X4 _209_ (
  .A(_119_),
  .Z(_120_)
);

NAND2_X1 _210_ (
  .A1(_118_),
  .A2(_120_),
  .ZN(_121_)
);

NAND2_X1 _211_ (
  .A1(_112_),
  .A2(_184_),
  .ZN(_122_)
);

INV_X1 _212_ (
  .A(_178_),
  .ZN(_123_)
);

NAND2_X1 _213_ (
  .A1(_123_),
  .A2(_106_),
  .ZN(_124_)
);

NAND3_X1 _214_ (
  .A1(_122_),
  .A2(_124_),
  .A3(_110_),
  .ZN(_125_)
);

INV_X1 _215_ (
  .A(_119_),
  .ZN(_126_)
);

BUF_X4 _216_ (
  .A(_126_),
  .Z(_127_)
);

BUF_X16 _217_ (
  .A(_116_),
  .Z(_128_)
);

NAND2_X1 _218_ (
  .A1(_128_),
  .A2(x[1]),
  .ZN(_129_)
);

NAND3_X1 _219_ (
  .A1(_125_),
  .A2(_127_),
  .A3(_129_),
  .ZN(_130_)
);

BUF_X2 _220_ (
  .A(y[2]),
  .Z(_131_)
);

BUF_X2 _221_ (
  .A(_131_),
  .Z(_132_)
);

NAND3_X1 _222_ (
  .A1(_121_),
  .A2(_130_),
  .A3(_132_),
  .ZN(_133_)
);

NAND2_X4 _223_ (
  .A1(_112_),
  .A2(_176_),
  .ZN(_134_)
);

INV_X1 _224_ (
  .A(_186_),
  .ZN(_135_)
);

NAND2_X1 _225_ (
  .A1(_135_),
  .A2(_106_),
  .ZN(_136_)
);

NAND2_X1 _226_ (
  .A1(_134_),
  .A2(_136_),
  .ZN(_137_)
);

NAND2_X2 _227_ (
  .A1(_137_),
  .A2(_110_),
  .ZN(_138_)
);

NAND3_X1 _228_ (
  .A1(_105_),
  .A2(_128_),
  .A3(_107_),
  .ZN(_139_)
);

NAND2_X1 _229_ (
  .A1(_138_),
  .A2(_139_),
  .ZN(_140_)
);

NAND2_X1 _230_ (
  .A1(_140_),
  .A2(_127_),
  .ZN(_141_)
);

INV_X1 _231_ (
  .A(_182_),
  .ZN(_142_)
);

NAND2_X1 _232_ (
  .A1(_103_),
  .A2(_142_),
  .ZN(_143_)
);

NAND2_X4 _233_ (
  .A1(_106_),
  .A2(_180_),
  .ZN(_144_)
);

NAND3_X1 _234_ (
  .A1(_143_),
  .A2(_128_),
  .A3(_144_),
  .ZN(_145_)
);

NAND2_X1 _235_ (
  .A1(_173_),
  .A2(_109_),
  .ZN(_146_)
);

NAND2_X1 _236_ (
  .A1(_146_),
  .A2(_119_),
  .ZN(_147_)
);

INV_X1 _237_ (
  .A(_147_),
  .ZN(_148_)
);

NAND2_X1 _238_ (
  .A1(_145_),
  .A2(_148_),
  .ZN(_149_)
);

INV_X1 _239_ (
  .A(_131_),
  .ZN(_150_)
);

NAND3_X1 _240_ (
  .A1(_141_),
  .A2(_149_),
  .A3(_150_),
  .ZN(_151_)
);

BUF_X4 _241_ (
  .A(ena),
  .Z(_152_)
);

NAND3_X1 _242_ (
  .A1(_133_),
  .A2(_151_),
  .A3(_152_),
  .ZN(_153_)
);

INV_X2 _243_ (
  .A(_152_),
  .ZN(_154_)
);

NAND2_X1 _244_ (
  .A1(_154_),
  .A2(\coef[21] ),
  .ZN(_155_)
);

NAND2_X1 _245_ (
  .A1(_153_),
  .A2(_155_),
  .ZN(_000_)
);

NAND2_X1 _246_ (
  .A1(_113_),
  .A2(_115_),
  .ZN(_156_)
);

NAND2_X1 _247_ (
  .A1(_156_),
  .A2(_110_),
  .ZN(_157_)
);

NAND3_X1 _248_ (
  .A1(_157_),
  .A2(_145_),
  .A3(_126_),
  .ZN(_158_)
);

AOI21_X1 _249_ (
  .A(_131_),
  .B1(_173_),
  .B2(_119_),
  .ZN(_159_)
);

AOI21_X1 _250_ (
  .A(_154_),
  .B1(_158_),
  .B2(_159_),
  .ZN(_160_)
);

NAND3_X1 _251_ (
  .A1(_134_),
  .A2(_136_),
  .A3(_128_),
  .ZN(_161_)
);

NAND3_X1 _252_ (
  .A1(_125_),
  .A2(_161_),
  .A3(_120_),
  .ZN(_162_)
);

NAND2_X1 _253_ (
  .A1(_127_),
  .A2(x[1]),
  .ZN(_009_)
);

NAND3_X1 _254_ (
  .A1(_162_),
  .A2(_132_),
  .A3(_009_),
  .ZN(_010_)
);

NAND2_X1 _255_ (
  .A1(_160_),
  .A2(_010_),
  .ZN(_011_)
);

INV_X1 _256_ (
  .A(\coef[23] ),
  .ZN(_012_)
);

OAI21_X1 _257_ (
  .A(_011_),
  .B1(_152_),
  .B2(_012_),
  .ZN(_001_)
);

NOR2_X1 _258_ (
  .A1(_152_),
  .A2(\coef[24] ),
  .ZN(_013_)
);

INV_X1 _259_ (
  .A(_184_),
  .ZN(_014_)
);

NAND2_X2 _260_ (
  .A1(_112_),
  .A2(_014_),
  .ZN(_015_)
);

NAND2_X1 _261_ (
  .A1(_106_),
  .A2(_178_),
  .ZN(_016_)
);

NAND3_X2 _262_ (
  .A1(_015_),
  .A2(_116_),
  .A3(_016_),
  .ZN(_017_)
);

AOI21_X1 _263_ (
  .A(_132_),
  .B1(_017_),
  .B2(_148_),
  .ZN(_018_)
);

NAND2_X1 _264_ (
  .A1(_112_),
  .A2(_178_),
  .ZN(_019_)
);

NAND2_X1 _265_ (
  .A1(_014_),
  .A2(_106_),
  .ZN(_020_)
);

NAND3_X1 _266_ (
  .A1(_019_),
  .A2(_020_),
  .A3(_128_),
  .ZN(_021_)
);

NAND2_X1 _267_ (
  .A1(_112_),
  .A2(_109_),
  .ZN(_022_)
);

NAND3_X1 _268_ (
  .A1(_021_),
  .A2(_127_),
  .A3(_022_),
  .ZN(_023_)
);

AOI21_X1 _269_ (
  .A(_154_),
  .B1(_018_),
  .B2(_023_),
  .ZN(_024_)
);

NAND2_X1 _270_ (
  .A1(_143_),
  .A2(_144_),
  .ZN(_025_)
);

NAND2_X2 _271_ (
  .A1(_025_),
  .A2(_109_),
  .ZN(_026_)
);

NAND3_X1 _272_ (
  .A1(_026_),
  .A2(_127_),
  .A3(_129_),
  .ZN(_027_)
);

INV_X1 _273_ (
  .A(_180_),
  .ZN(_028_)
);

NAND2_X1 _274_ (
  .A1(_112_),
  .A2(_028_),
  .ZN(_029_)
);

NAND2_X1 _275_ (
  .A1(_106_),
  .A2(_182_),
  .ZN(_030_)
);

NAND3_X1 _276_ (
  .A1(_029_),
  .A2(_110_),
  .A3(_030_),
  .ZN(_031_)
);

NOR2_X1 _277_ (
  .A1(_112_),
  .A2(_109_),
  .ZN(_032_)
);

INV_X1 _278_ (
  .A(_032_),
  .ZN(_033_)
);

NAND3_X1 _279_ (
  .A1(_031_),
  .A2(_120_),
  .A3(_033_),
  .ZN(_034_)
);

NAND3_X1 _280_ (
  .A1(_027_),
  .A2(_034_),
  .A3(_132_),
  .ZN(_035_)
);

AOI21_X1 _281_ (
  .A(_013_),
  .B1(_024_),
  .B2(_035_),
  .ZN(_002_)
);

NAND3_X1 _282_ (
  .A1(_111_),
  .A2(_120_),
  .A3(_033_),
  .ZN(_036_)
);

AOI21_X2 _283_ (
  .A(_119_),
  .B1(_128_),
  .B2(x[0]),
  .ZN(_037_)
);

AOI21_X1 _284_ (
  .A(_131_),
  .B1(_037_),
  .B2(_146_),
  .ZN(_038_)
);

AOI21_X1 _285_ (
  .A(_154_),
  .B1(_036_),
  .B2(_038_),
  .ZN(_039_)
);

NAND3_X1 _286_ (
  .A1(_139_),
  .A2(_126_),
  .A3(_022_),
  .ZN(_040_)
);

NAND2_X1 _287_ (
  .A1(_172_),
  .A2(_110_),
  .ZN(_041_)
);

NAND3_X1 _288_ (
  .A1(_129_),
  .A2(_041_),
  .A3(_119_),
  .ZN(_042_)
);

NAND3_X1 _289_ (
  .A1(_040_),
  .A2(_132_),
  .A3(_042_),
  .ZN(_043_)
);

NAND2_X1 _290_ (
  .A1(_039_),
  .A2(_043_),
  .ZN(_044_)
);

INV_X1 _291_ (
  .A(\coef[10] ),
  .ZN(_045_)
);

OAI21_X1 _292_ (
  .A(_044_),
  .B1(_152_),
  .B2(_045_),
  .ZN(_003_)
);

NAND2_X1 _293_ (
  .A1(_108_),
  .A2(_128_),
  .ZN(_046_)
);

NAND3_X1 _294_ (
  .A1(_157_),
  .A2(_046_),
  .A3(_127_),
  .ZN(_047_)
);

NAND2_X1 _295_ (
  .A1(_138_),
  .A2(_129_),
  .ZN(_048_)
);

NAND2_X1 _296_ (
  .A1(_048_),
  .A2(_120_),
  .ZN(_049_)
);

NAND3_X1 _297_ (
  .A1(_047_),
  .A2(_049_),
  .A3(_132_),
  .ZN(_050_)
);

NAND2_X1 _298_ (
  .A1(_117_),
  .A2(_146_),
  .ZN(_051_)
);

NAND2_X1 _299_ (
  .A1(_051_),
  .A2(_127_),
  .ZN(_052_)
);

NAND3_X1 _300_ (
  .A1(_105_),
  .A2(_110_),
  .A3(_107_),
  .ZN(_053_)
);

NAND3_X1 _301_ (
  .A1(_161_),
  .A2(_053_),
  .A3(_120_),
  .ZN(_054_)
);

NAND3_X1 _302_ (
  .A1(_052_),
  .A2(_054_),
  .A3(_150_),
  .ZN(_055_)
);

NAND3_X1 _303_ (
  .A1(_050_),
  .A2(_055_),
  .A3(_152_),
  .ZN(_056_)
);

NAND2_X1 _304_ (
  .A1(_154_),
  .A2(\coef[26] ),
  .ZN(_057_)
);

NAND2_X1 _305_ (
  .A1(_056_),
  .A2(_057_),
  .ZN(_004_)
);

NOR2_X1 _306_ (
  .A1(_152_),
  .A2(\coef[13] ),
  .ZN(_058_)
);

NAND3_X1 _307_ (
  .A1(_019_),
  .A2(_020_),
  .A3(_110_),
  .ZN(_059_)
);

AOI21_X1 _308_ (
  .A(_132_),
  .B1(_059_),
  .B2(_037_),
  .ZN(_060_)
);

NAND2_X1 _309_ (
  .A1(_112_),
  .A2(_114_),
  .ZN(_061_)
);

NAND2_X1 _310_ (
  .A1(_106_),
  .A2(_174_),
  .ZN(_062_)
);

NAND3_X1 _311_ (
  .A1(_061_),
  .A2(_128_),
  .A3(_062_),
  .ZN(_063_)
);

NAND2_X1 _312_ (
  .A1(_022_),
  .A2(_119_),
  .ZN(_064_)
);

INV_X1 _313_ (
  .A(_064_),
  .ZN(_065_)
);

NAND2_X1 _314_ (
  .A1(_063_),
  .A2(_065_),
  .ZN(_066_)
);

AOI21_X1 _315_ (
  .A(_154_),
  .B1(_060_),
  .B2(_066_),
  .ZN(_067_)
);

NAND3_X1 _316_ (
  .A1(_029_),
  .A2(_128_),
  .A3(_030_),
  .ZN(_068_)
);

NAND3_X1 _317_ (
  .A1(_068_),
  .A2(_120_),
  .A3(_041_),
  .ZN(_069_)
);

NAND2_X1 _318_ (
  .A1(_112_),
  .A2(_186_),
  .ZN(_070_)
);

INV_X1 _319_ (
  .A(_176_),
  .ZN(_071_)
);

NAND2_X1 _320_ (
  .A1(_071_),
  .A2(_106_),
  .ZN(_072_)
);

NAND3_X1 _321_ (
  .A1(_070_),
  .A2(_072_),
  .A3(_110_),
  .ZN(_073_)
);

NOR2_X1 _322_ (
  .A1(_032_),
  .A2(_119_),
  .ZN(_074_)
);

NAND2_X1 _323_ (
  .A1(_073_),
  .A2(_074_),
  .ZN(_075_)
);

NAND3_X1 _324_ (
  .A1(_069_),
  .A2(_132_),
  .A3(_075_),
  .ZN(_076_)
);

AOI21_X1 _325_ (
  .A(_058_),
  .B1(_067_),
  .B2(_076_),
  .ZN(_005_)
);

NAND3_X1 _326_ (
  .A1(_021_),
  .A2(_073_),
  .A3(_126_),
  .ZN(_077_)
);

NAND3_X1 _327_ (
  .A1(_138_),
  .A2(_017_),
  .A3(_119_),
  .ZN(_078_)
);

NAND3_X1 _328_ (
  .A1(_077_),
  .A2(_078_),
  .A3(_150_),
  .ZN(_079_)
);

NAND3_X1 _329_ (
  .A1(_026_),
  .A2(_117_),
  .A3(_126_),
  .ZN(_080_)
);

NAND3_X1 _330_ (
  .A1(_031_),
  .A2(_063_),
  .A3(_119_),
  .ZN(_081_)
);

NAND3_X1 _331_ (
  .A1(_080_),
  .A2(_081_),
  .A3(_132_),
  .ZN(_082_)
);

NAND2_X1 _332_ (
  .A1(_079_),
  .A2(_082_),
  .ZN(_083_)
);

NAND2_X1 _333_ (
  .A1(_083_),
  .A2(_152_),
  .ZN(_084_)
);

NAND2_X1 _334_ (
  .A1(_154_),
  .A2(\coef[28] ),
  .ZN(_085_)
);

NAND2_X2 _335_ (
  .A1(_084_),
  .A2(_085_),
  .ZN(_006_)
);

NOR2_X1 _336_ (
  .A1(_152_),
  .A2(\coef[29] ),
  .ZN(_086_)
);

AOI21_X1 _337_ (
  .A(_131_),
  .B1(_053_),
  .B2(_074_),
  .ZN(_087_)
);

NAND3_X1 _338_ (
  .A1(_061_),
  .A2(_110_),
  .A3(_062_),
  .ZN(_088_)
);

NAND3_X1 _339_ (
  .A1(_017_),
  .A2(_088_),
  .A3(_120_),
  .ZN(_089_)
);

AOI21_X1 _340_ (
  .A(_154_),
  .B1(_087_),
  .B2(_089_),
  .ZN(_090_)
);

AOI21_X1 _341_ (
  .A(_150_),
  .B1(_046_),
  .B2(_065_),
  .ZN(_091_)
);

NAND3_X1 _342_ (
  .A1(_070_),
  .A2(_072_),
  .A3(_128_),
  .ZN(_092_)
);

NAND3_X1 _343_ (
  .A1(_026_),
  .A2(_092_),
  .A3(_127_),
  .ZN(_093_)
);

NAND2_X1 _344_ (
  .A1(_091_),
  .A2(_093_),
  .ZN(_094_)
);

AOI21_X2 _345_ (
  .A(_086_),
  .B1(_090_),
  .B2(_094_),
  .ZN(_007_)
);

NOR2_X1 _346_ (
  .A1(_152_),
  .A2(\coef[30] ),
  .ZN(_095_)
);

NAND3_X1 _347_ (
  .A1(_026_),
  .A2(_017_),
  .A3(_127_),
  .ZN(_096_)
);

NAND2_X1 _348_ (
  .A1(_015_),
  .A2(_016_),
  .ZN(_097_)
);

AOI21_X1 _349_ (
  .A(_131_),
  .B1(_097_),
  .B2(_120_),
  .ZN(_098_)
);

AOI21_X1 _350_ (
  .A(_154_),
  .B1(_096_),
  .B2(_098_),
  .ZN(_099_)
);

NAND3_X1 _351_ (
  .A1(_026_),
  .A2(_017_),
  .A3(_120_),
  .ZN(_100_)
);

NAND3_X1 _352_ (
  .A1(_143_),
  .A2(_127_),
  .A3(_144_),
  .ZN(_101_)
);

NAND3_X1 _353_ (
  .A1(_100_),
  .A2(_132_),
  .A3(_101_),
  .ZN(_102_)
);

AOI21_X1 _354_ (
  .A(_095_),
  .B1(_099_),
  .B2(_102_),
  .ZN(_008_)
);

HA_X1 _355_ (
  .A(_172_),
  .B(_173_),
  .CO(_174_),
  .S(_175_)
);

HA_X1 _356_ (
  .A(_172_),
  .B(_173_),
  .CO(_176_),
  .S(_177_)
);

HA_X1 _357_ (
  .A(_172_),
  .B(x[1]),
  .CO(_178_),
  .S(_179_)
);

HA_X1 _358_ (
  .A(_172_),
  .B(x[1]),
  .CO(_180_),
  .S(_181_)
);

HA_X1 _359_ (
  .A(x[0]),
  .B(_173_),
  .CO(_182_),
  .S(_183_)
);

HA_X1 _360_ (
  .A(x[0]),
  .B(_173_),
  .CO(_184_),
  .S(_185_)
);

HA_X1 _361_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_186_),
  .S(_187_)
);

HA_X1 _362_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_188_),
  .S(_189_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_171_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_170_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_169_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_168_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_167_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_166_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_165_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_164_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_163_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$bfc28a02cfebf191b4a982c9147f38f65a3f3469\dctu

module \$paramod$c4f8cc56c0ef9356356d2a98d35862f209dd307b\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _177_ (
  .A(x[0]),
  .ZN(_159_)
);

INV_X1 _178_ (
  .A(x[1]),
  .ZN(_160_)
);

CLKBUF_X3 _179_ (
  .A(ena),
  .Z(_091_)
);

NOR2_X1 _180_ (
  .A1(\coef[21] ),
  .A2(_091_),
  .ZN(_092_)
);

INV_X2 _181_ (
  .A(_091_),
  .ZN(_093_)
);

INV_X2 _182_ (
  .A(x[2]),
  .ZN(_094_)
);

XNOR2_X2 _183_ (
  .A(_094_),
  .B(_162_),
  .ZN(_095_)
);

INV_X2 _184_ (
  .A(_095_),
  .ZN(_096_)
);

BUF_X4 _185_ (
  .A(y[0]),
  .Z(_097_)
);

BUF_X4 _186_ (
  .A(_097_),
  .Z(_098_)
);

NAND2_X1 _187_ (
  .A1(_096_),
  .A2(_098_),
  .ZN(_099_)
);

BUF_X2 _188_ (
  .A(y[1]),
  .Z(_100_)
);

BUF_X4 _189_ (
  .A(_100_),
  .Z(_101_)
);

BUF_X4 _190_ (
  .A(_101_),
  .Z(_102_)
);

BUF_X8 _191_ (
  .A(_094_),
  .Z(_103_)
);

INV_X1 _192_ (
  .A(_163_),
  .ZN(_104_)
);

NAND2_X4 _193_ (
  .A1(_103_),
  .A2(_104_),
  .ZN(_105_)
);

INV_X8 _194_ (
  .A(_097_),
  .ZN(_106_)
);

BUF_X8 _195_ (
  .A(_106_),
  .Z(_107_)
);

BUF_X4 _196_ (
  .A(x[2]),
  .Z(_108_)
);

NAND2_X2 _197_ (
  .A1(_108_),
  .A2(_173_),
  .ZN(_109_)
);

NAND3_X1 _198_ (
  .A1(_105_),
  .A2(_107_),
  .A3(_109_),
  .ZN(_110_)
);

NAND3_X1 _199_ (
  .A1(_099_),
  .A2(_102_),
  .A3(_110_),
  .ZN(_111_)
);

CLKBUF_X3 _200_ (
  .A(y[2]),
  .Z(_112_)
);

INV_X1 _201_ (
  .A(_171_),
  .ZN(_113_)
);

NAND2_X4 _202_ (
  .A1(_103_),
  .A2(_113_),
  .ZN(_114_)
);

NAND2_X1 _203_ (
  .A1(_108_),
  .A2(_165_),
  .ZN(_115_)
);

NAND3_X2 _204_ (
  .A1(_114_),
  .A2(_097_),
  .A3(_115_),
  .ZN(_116_)
);

AOI21_X2 _205_ (
  .A(_101_),
  .B1(_106_),
  .B2(x[1]),
  .ZN(_117_)
);

AOI21_X1 _206_ (
  .A(_112_),
  .B1(_116_),
  .B2(_117_),
  .ZN(_118_)
);

AOI21_X1 _207_ (
  .A(_093_),
  .B1(_111_),
  .B2(_118_),
  .ZN(_119_)
);

NAND2_X2 _208_ (
  .A1(_095_),
  .A2(_106_),
  .ZN(_120_)
);

INV_X1 _209_ (
  .A(_100_),
  .ZN(_121_)
);

NAND2_X4 _210_ (
  .A1(_103_),
  .A2(_161_),
  .ZN(_122_)
);

INV_X1 _211_ (
  .A(_175_),
  .ZN(_123_)
);

NAND2_X2 _212_ (
  .A1(_123_),
  .A2(_108_),
  .ZN(_124_)
);

NAND3_X1 _213_ (
  .A1(_122_),
  .A2(_124_),
  .A3(_098_),
  .ZN(_125_)
);

NAND3_X1 _214_ (
  .A1(_120_),
  .A2(_121_),
  .A3(_125_),
  .ZN(_126_)
);

INV_X2 _215_ (
  .A(_112_),
  .ZN(_127_)
);

NAND2_X2 _216_ (
  .A1(_103_),
  .A2(_169_),
  .ZN(_128_)
);

INV_X1 _217_ (
  .A(_167_),
  .ZN(_129_)
);

NAND2_X1 _218_ (
  .A1(_129_),
  .A2(_108_),
  .ZN(_130_)
);

NAND3_X2 _219_ (
  .A1(_128_),
  .A2(_130_),
  .A3(_106_),
  .ZN(_131_)
);

OAI21_X1 _220_ (
  .A(_100_),
  .B1(_106_),
  .B2(x[1]),
  .ZN(_132_)
);

INV_X1 _221_ (
  .A(_132_),
  .ZN(_133_)
);

AOI21_X1 _222_ (
  .A(_127_),
  .B1(_131_),
  .B2(_133_),
  .ZN(_134_)
);

NAND2_X1 _223_ (
  .A1(_126_),
  .A2(_134_),
  .ZN(_135_)
);

AOI21_X2 _224_ (
  .A(_092_),
  .B1(_119_),
  .B2(_135_),
  .ZN(_000_)
);

NOR2_X1 _225_ (
  .A1(_091_),
  .A2(\coef[23] ),
  .ZN(_136_)
);

AOI21_X1 _226_ (
  .A(_112_),
  .B1(_096_),
  .B2(_102_),
  .ZN(_137_)
);

NAND3_X1 _227_ (
  .A1(_128_),
  .A2(_130_),
  .A3(_098_),
  .ZN(_138_)
);

NAND3_X1 _228_ (
  .A1(_138_),
  .A2(_110_),
  .A3(_121_),
  .ZN(_139_)
);

AOI21_X1 _229_ (
  .A(_093_),
  .B1(_137_),
  .B2(_139_),
  .ZN(_140_)
);

NAND3_X1 _230_ (
  .A1(_114_),
  .A2(_107_),
  .A3(_115_),
  .ZN(_141_)
);

NAND3_X1 _231_ (
  .A1(_125_),
  .A2(_141_),
  .A3(_102_),
  .ZN(_142_)
);

AOI21_X1 _232_ (
  .A(_127_),
  .B1(_095_),
  .B2(_121_),
  .ZN(_143_)
);

NAND2_X1 _233_ (
  .A1(_142_),
  .A2(_143_),
  .ZN(_144_)
);

AOI21_X1 _234_ (
  .A(_136_),
  .B1(_140_),
  .B2(_144_),
  .ZN(_001_)
);

NOR2_X1 _235_ (
  .A1(_091_),
  .A2(\coef[24] ),
  .ZN(_145_)
);

NAND2_X2 _236_ (
  .A1(_096_),
  .A2(_107_),
  .ZN(_146_)
);

NAND3_X4 _237_ (
  .A1(_105_),
  .A2(_097_),
  .A3(_109_),
  .ZN(_147_)
);

NAND3_X1 _238_ (
  .A1(_146_),
  .A2(_121_),
  .A3(_147_),
  .ZN(_148_)
);

NAND2_X2 _239_ (
  .A1(_103_),
  .A2(_123_),
  .ZN(_149_)
);

NAND2_X1 _240_ (
  .A1(_108_),
  .A2(_161_),
  .ZN(_009_)
);

NAND3_X2 _241_ (
  .A1(_149_),
  .A2(_098_),
  .A3(_009_),
  .ZN(_010_)
);

NAND2_X1 _242_ (
  .A1(_106_),
  .A2(x[0]),
  .ZN(_011_)
);

NAND2_X1 _243_ (
  .A1(_011_),
  .A2(_101_),
  .ZN(_012_)
);

INV_X1 _244_ (
  .A(_012_),
  .ZN(_013_)
);

AOI21_X1 _245_ (
  .A(_127_),
  .B1(_010_),
  .B2(_013_),
  .ZN(_014_)
);

AOI21_X1 _246_ (
  .A(_093_),
  .B1(_148_),
  .B2(_014_),
  .ZN(_015_)
);

NAND3_X4 _247_ (
  .A1(_122_),
  .A2(_124_),
  .A3(_106_),
  .ZN(_016_)
);

AND2_X4 _248_ (
  .A1(_016_),
  .A2(_101_),
  .ZN(_017_)
);

NAND2_X2 _249_ (
  .A1(_095_),
  .A2(_098_),
  .ZN(_018_)
);

NAND2_X2 _250_ (
  .A1(_017_),
  .A2(_018_),
  .ZN(_019_)
);

NAND2_X2 _251_ (
  .A1(_103_),
  .A2(_173_),
  .ZN(_020_)
);

NAND2_X1 _252_ (
  .A1(_104_),
  .A2(_108_),
  .ZN(_021_)
);

NAND3_X1 _253_ (
  .A1(_020_),
  .A2(_021_),
  .A3(_106_),
  .ZN(_022_)
);

NAND2_X1 _254_ (
  .A1(_159_),
  .A2(_097_),
  .ZN(_023_)
);

NAND3_X1 _255_ (
  .A1(_022_),
  .A2(_121_),
  .A3(_023_),
  .ZN(_024_)
);

NAND3_X2 _256_ (
  .A1(_019_),
  .A2(_127_),
  .A3(_024_),
  .ZN(_025_)
);

AOI21_X2 _257_ (
  .A(_145_),
  .B1(_015_),
  .B2(_025_),
  .ZN(_002_)
);

NAND2_X1 _258_ (
  .A1(_103_),
  .A2(_107_),
  .ZN(_026_)
);

NAND3_X1 _259_ (
  .A1(_018_),
  .A2(_121_),
  .A3(_026_),
  .ZN(_027_)
);

AOI21_X1 _260_ (
  .A(_112_),
  .B1(_133_),
  .B2(_011_),
  .ZN(_028_)
);

AOI21_X1 _261_ (
  .A(_093_),
  .B1(_027_),
  .B2(_028_),
  .ZN(_029_)
);

OAI21_X1 _262_ (
  .A(_120_),
  .B1(_108_),
  .B2(_107_),
  .ZN(_030_)
);

NAND2_X1 _263_ (
  .A1(_030_),
  .A2(_102_),
  .ZN(_031_)
);

AOI21_X1 _264_ (
  .A(_127_),
  .B1(_117_),
  .B2(_023_),
  .ZN(_032_)
);

NAND2_X1 _265_ (
  .A1(_031_),
  .A2(_032_),
  .ZN(_033_)
);

NAND2_X1 _266_ (
  .A1(_029_),
  .A2(_033_),
  .ZN(_034_)
);

NAND2_X1 _267_ (
  .A1(_093_),
  .A2(\coef[10] ),
  .ZN(_035_)
);

NAND2_X1 _268_ (
  .A1(_034_),
  .A2(_035_),
  .ZN(_003_)
);

NOR2_X1 _269_ (
  .A1(_091_),
  .A2(\coef[26] ),
  .ZN(_036_)
);

NAND3_X1 _270_ (
  .A1(_018_),
  .A2(_121_),
  .A3(_131_),
  .ZN(_037_)
);

AOI21_X1 _271_ (
  .A(_112_),
  .B1(_141_),
  .B2(_133_),
  .ZN(_038_)
);

AOI21_X1 _272_ (
  .A(_093_),
  .B1(_037_),
  .B2(_038_),
  .ZN(_039_)
);

NAND3_X1 _273_ (
  .A1(_146_),
  .A2(_102_),
  .A3(_116_),
  .ZN(_040_)
);

AOI21_X1 _274_ (
  .A(_127_),
  .B1(_138_),
  .B2(_117_),
  .ZN(_041_)
);

NAND2_X1 _275_ (
  .A1(_040_),
  .A2(_041_),
  .ZN(_042_)
);

AOI21_X2 _276_ (
  .A(_036_),
  .B1(_039_),
  .B2(_042_),
  .ZN(_004_)
);

NOR2_X1 _277_ (
  .A1(_091_),
  .A2(\coef[13] ),
  .ZN(_043_)
);

NAND3_X1 _278_ (
  .A1(_020_),
  .A2(_021_),
  .A3(_098_),
  .ZN(_044_)
);

AOI21_X1 _279_ (
  .A(_101_),
  .B1(_107_),
  .B2(_103_),
  .ZN(_045_)
);

AOI21_X1 _280_ (
  .A(_112_),
  .B1(_044_),
  .B2(_045_),
  .ZN(_046_)
);

NAND2_X2 _281_ (
  .A1(_103_),
  .A2(_165_),
  .ZN(_047_)
);

NAND2_X1 _282_ (
  .A1(_113_),
  .A2(_108_),
  .ZN(_048_)
);

NAND3_X1 _283_ (
  .A1(_047_),
  .A2(_048_),
  .A3(_106_),
  .ZN(_049_)
);

NAND3_X1 _284_ (
  .A1(_049_),
  .A2(_102_),
  .A3(_023_),
  .ZN(_050_)
);

AOI21_X1 _285_ (
  .A(_093_),
  .B1(_046_),
  .B2(_050_),
  .ZN(_051_)
);

NAND2_X2 _286_ (
  .A1(_103_),
  .A2(_129_),
  .ZN(_052_)
);

NAND2_X1 _287_ (
  .A1(_108_),
  .A2(_169_),
  .ZN(_053_)
);

NAND3_X2 _288_ (
  .A1(_052_),
  .A2(_098_),
  .A3(_053_),
  .ZN(_054_)
);

AOI21_X4 _289_ (
  .A(_101_),
  .B1(_107_),
  .B2(x[0]),
  .ZN(_055_)
);

AOI21_X1 _290_ (
  .A(_127_),
  .B1(_054_),
  .B2(_055_),
  .ZN(_056_)
);

NAND3_X1 _291_ (
  .A1(_149_),
  .A2(_107_),
  .A3(_009_),
  .ZN(_057_)
);

NAND2_X1 _292_ (
  .A1(_108_),
  .A2(_098_),
  .ZN(_058_)
);

NAND3_X1 _293_ (
  .A1(_057_),
  .A2(_102_),
  .A3(_058_),
  .ZN(_059_)
);

NAND2_X1 _294_ (
  .A1(_056_),
  .A2(_059_),
  .ZN(_060_)
);

AOI21_X1 _295_ (
  .A(_043_),
  .B1(_051_),
  .B2(_060_),
  .ZN(_005_)
);

NAND3_X1 _296_ (
  .A1(_022_),
  .A2(_054_),
  .A3(_121_),
  .ZN(_061_)
);

NAND3_X1 _297_ (
  .A1(_016_),
  .A2(_116_),
  .A3(_101_),
  .ZN(_062_)
);

NAND3_X1 _298_ (
  .A1(_061_),
  .A2(_062_),
  .A3(_127_),
  .ZN(_063_)
);

NAND3_X1 _299_ (
  .A1(_131_),
  .A2(_147_),
  .A3(_121_),
  .ZN(_064_)
);

NAND3_X1 _300_ (
  .A1(_049_),
  .A2(_010_),
  .A3(_101_),
  .ZN(_065_)
);

NAND3_X1 _301_ (
  .A1(_064_),
  .A2(_065_),
  .A3(_112_),
  .ZN(_066_)
);

NAND2_X1 _302_ (
  .A1(_063_),
  .A2(_066_),
  .ZN(_067_)
);

NAND2_X1 _303_ (
  .A1(_067_),
  .A2(_091_),
  .ZN(_068_)
);

NAND2_X1 _304_ (
  .A1(_093_),
  .A2(\coef[28] ),
  .ZN(_069_)
);

NAND2_X1 _305_ (
  .A1(_068_),
  .A2(_069_),
  .ZN(_006_)
);

NAND2_X1 _306_ (
  .A1(_093_),
  .A2(\coef[29] ),
  .ZN(_070_)
);

NAND3_X1 _307_ (
  .A1(_052_),
  .A2(_107_),
  .A3(_053_),
  .ZN(_071_)
);

AOI21_X1 _308_ (
  .A(_102_),
  .B1(_147_),
  .B2(_071_),
  .ZN(_072_)
);

OAI21_X1 _309_ (
  .A(_023_),
  .B1(_098_),
  .B2(x[1]),
  .ZN(_073_)
);

NAND2_X1 _310_ (
  .A1(_073_),
  .A2(_102_),
  .ZN(_074_)
);

NAND2_X1 _311_ (
  .A1(_074_),
  .A2(_112_),
  .ZN(_075_)
);

OAI21_X1 _312_ (
  .A(_091_),
  .B1(_072_),
  .B2(_075_),
  .ZN(_076_)
);

NAND3_X1 _313_ (
  .A1(_047_),
  .A2(_048_),
  .A3(_098_),
  .ZN(_077_)
);

NAND3_X1 _314_ (
  .A1(_016_),
  .A2(_077_),
  .A3(_102_),
  .ZN(_078_)
);

OAI21_X1 _315_ (
  .A(_055_),
  .B1(_107_),
  .B2(_160_),
  .ZN(_079_)
);

AOI21_X1 _316_ (
  .A(_112_),
  .B1(_078_),
  .B2(_079_),
  .ZN(_080_)
);

OAI21_X2 _317_ (
  .A(_070_),
  .B1(_076_),
  .B2(_080_),
  .ZN(_007_)
);

AND2_X1 _318_ (
  .A1(_147_),
  .A2(_112_),
  .ZN(_081_)
);

AOI21_X1 _319_ (
  .A(_101_),
  .B1(_105_),
  .B2(_109_),
  .ZN(_082_)
);

OAI21_X2 _320_ (
  .A(_081_),
  .B1(_017_),
  .B2(_082_),
  .ZN(_083_)
);

NAND2_X1 _321_ (
  .A1(_147_),
  .A2(_121_),
  .ZN(_084_)
);

NAND2_X1 _322_ (
  .A1(_122_),
  .A2(_124_),
  .ZN(_085_)
);

NAND2_X1 _323_ (
  .A1(_085_),
  .A2(_101_),
  .ZN(_086_)
);

NAND2_X1 _324_ (
  .A1(_084_),
  .A2(_086_),
  .ZN(_087_)
);

NAND3_X1 _325_ (
  .A1(_087_),
  .A2(_127_),
  .A3(_016_),
  .ZN(_088_)
);

NAND3_X1 _326_ (
  .A1(_083_),
  .A2(_088_),
  .A3(_091_),
  .ZN(_089_)
);

NAND2_X1 _327_ (
  .A1(_093_),
  .A2(\coef[30] ),
  .ZN(_090_)
);

NAND2_X1 _328_ (
  .A1(_089_),
  .A2(_090_),
  .ZN(_008_)
);

HA_X1 _329_ (
  .A(_159_),
  .B(_160_),
  .CO(_161_),
  .S(_162_)
);

HA_X1 _330_ (
  .A(_159_),
  .B(_160_),
  .CO(_163_),
  .S(_164_)
);

HA_X1 _331_ (
  .A(_159_),
  .B(x[1]),
  .CO(_165_),
  .S(_166_)
);

HA_X1 _332_ (
  .A(_159_),
  .B(x[1]),
  .CO(_167_),
  .S(_168_)
);

HA_X1 _333_ (
  .A(x[0]),
  .B(_160_),
  .CO(_169_),
  .S(_170_)
);

HA_X1 _334_ (
  .A(x[0]),
  .B(_160_),
  .CO(_171_),
  .S(_172_)
);

HA_X1 _335_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _336_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_175_),
  .S(_176_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_158_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_157_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_156_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_155_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_154_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_153_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_152_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_151_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_150_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$c4f8cc56c0ef9356356d2a98d35862f209dd307b\dctu

module \$paramod$c50cce30a10e9eb82ea37b86647b55ab680286c8\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire \coef[10] ;
wire \coef[11] ;
wire \coef[13] ;
wire \coef[15] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

BUF_X4 _30_ (
  .A(x[2]),
  .Z(_04_)
);

INV_X4 _31_ (
  .A(_04_),
  .ZN(_05_)
);

NAND2_X2 _32_ (
  .A1(_05_),
  .A2(x[0]),
  .ZN(_06_)
);

INV_X1 _33_ (
  .A(x[0]),
  .ZN(_07_)
);

NAND2_X1 _34_ (
  .A1(_07_),
  .A2(_04_),
  .ZN(_08_)
);

BUF_X4 _35_ (
  .A(ena),
  .Z(_09_)
);

NAND3_X1 _36_ (
  .A1(_06_),
  .A2(_08_),
  .A3(_09_),
  .ZN(_10_)
);

INV_X2 _37_ (
  .A(_09_),
  .ZN(_11_)
);

NAND2_X1 _38_ (
  .A1(_11_),
  .A2(\coef[11] ),
  .ZN(_12_)
);

NAND2_X1 _39_ (
  .A1(_10_),
  .A2(_12_),
  .ZN(_00_)
);

INV_X1 _40_ (
  .A(x[1]),
  .ZN(_13_)
);

NAND2_X1 _41_ (
  .A1(_13_),
  .A2(_04_),
  .ZN(_14_)
);

NAND2_X2 _42_ (
  .A1(_05_),
  .A2(x[1]),
  .ZN(_15_)
);

NAND3_X2 _43_ (
  .A1(_14_),
  .A2(_15_),
  .A3(_09_),
  .ZN(_16_)
);

NAND2_X1 _44_ (
  .A1(_11_),
  .A2(\coef[13] ),
  .ZN(_17_)
);

NAND2_X2 _45_ (
  .A1(_16_),
  .A2(_17_),
  .ZN(_01_)
);

NAND2_X1 _46_ (
  .A1(_11_),
  .A2(\coef[10] ),
  .ZN(_18_)
);

NAND2_X1 _47_ (
  .A1(_04_),
  .A2(x[1]),
  .ZN(_19_)
);

NAND2_X1 _48_ (
  .A1(_19_),
  .A2(_09_),
  .ZN(_20_)
);

NOR2_X1 _49_ (
  .A1(_04_),
  .A2(x[1]),
  .ZN(_21_)
);

OAI21_X2 _50_ (
  .A(_18_),
  .B1(_20_),
  .B2(_21_),
  .ZN(_02_)
);

NAND2_X1 _51_ (
  .A1(_11_),
  .A2(\coef[15] ),
  .ZN(_22_)
);

NAND2_X1 _52_ (
  .A1(_04_),
  .A2(x[0]),
  .ZN(_23_)
);

NAND2_X1 _53_ (
  .A1(_23_),
  .A2(_09_),
  .ZN(_24_)
);

NOR2_X1 _54_ (
  .A1(_04_),
  .A2(x[0]),
  .ZN(_25_)
);

OAI21_X2 _55_ (
  .A(_22_),
  .B1(_24_),
  .B2(_25_),
  .ZN(_03_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[11] ),
  .QN(_29_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_01_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_28_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_02_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_27_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_03_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_26_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[15] , \coef[15] , \coef[10] , \coef[13] , \coef[10] , \coef[15] , \coef[15] , \coef[11] , \coef[10] , \coef[11] , \coef[15] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$c50cce30a10e9eb82ea37b86647b55ab680286c8\dctu

module \$paramod$ca051f171e86125a3bcf4bd090f5be774b98c04e\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _184_ (
  .A(x[1]),
  .ZN(_167_)
);

INV_X1 _185_ (
  .A(x[0]),
  .ZN(_166_)
);

BUF_X2 _186_ (
  .A(y[2]),
  .Z(_097_)
);

INV_X1 _187_ (
  .A(_097_),
  .ZN(_098_)
);

BUF_X8 _188_ (
  .A(x[2]),
  .Z(_099_)
);

INV_X8 _189_ (
  .A(_099_),
  .ZN(_100_)
);

INV_X1 _190_ (
  .A(_174_),
  .ZN(_101_)
);

NAND2_X1 _191_ (
  .A1(_100_),
  .A2(_101_),
  .ZN(_102_)
);

BUF_X8 _192_ (
  .A(y[0]),
  .Z(_103_)
);

BUF_X16 _193_ (
  .A(_099_),
  .Z(_104_)
);

NAND2_X4 _194_ (
  .A1(_104_),
  .A2(_176_),
  .ZN(_105_)
);

NAND3_X2 _195_ (
  .A1(_102_),
  .A2(_103_),
  .A3(_105_),
  .ZN(_106_)
);

BUF_X4 _196_ (
  .A(y[1]),
  .Z(_107_)
);

BUF_X2 _197_ (
  .A(_107_),
  .Z(_108_)
);

INV_X4 _198_ (
  .A(y[0]),
  .ZN(_109_)
);

NAND2_X2 _199_ (
  .A1(_109_),
  .A2(_104_),
  .ZN(_110_)
);

NAND3_X1 _200_ (
  .A1(_106_),
  .A2(_108_),
  .A3(_110_),
  .ZN(_111_)
);

INV_X1 _201_ (
  .A(_111_),
  .ZN(_112_)
);

INV_X1 _202_ (
  .A(_180_),
  .ZN(_113_)
);

NAND2_X1 _203_ (
  .A1(_100_),
  .A2(_113_),
  .ZN(_114_)
);

BUF_X8 _204_ (
  .A(_109_),
  .Z(_115_)
);

NAND2_X4 _205_ (
  .A1(_104_),
  .A2(_170_),
  .ZN(_116_)
);

NAND3_X2 _206_ (
  .A1(_114_),
  .A2(_115_),
  .A3(_116_),
  .ZN(_117_)
);

NAND2_X1 _207_ (
  .A1(_166_),
  .A2(_103_),
  .ZN(_118_)
);

AOI21_X1 _208_ (
  .A(_108_),
  .B1(_117_),
  .B2(_118_),
  .ZN(_119_)
);

OAI21_X1 _209_ (
  .A(_098_),
  .B1(_112_),
  .B2(_119_),
  .ZN(_120_)
);

BUF_X2 _210_ (
  .A(ena),
  .Z(_121_)
);

INV_X2 _211_ (
  .A(_121_),
  .ZN(_122_)
);

INV_X1 _212_ (
  .A(_182_),
  .ZN(_123_)
);

NAND2_X2 _213_ (
  .A1(_100_),
  .A2(_123_),
  .ZN(_124_)
);

NAND2_X4 _214_ (
  .A1(_104_),
  .A2(_168_),
  .ZN(_125_)
);

NAND2_X2 _215_ (
  .A1(_124_),
  .A2(_125_),
  .ZN(_126_)
);

BUF_X16 _216_ (
  .A(_103_),
  .Z(_127_)
);

NAND2_X1 _217_ (
  .A1(_126_),
  .A2(_127_),
  .ZN(_128_)
);

NAND2_X2 _218_ (
  .A1(_109_),
  .A2(x[0]),
  .ZN(_129_)
);

NAND2_X1 _219_ (
  .A1(_129_),
  .A2(_107_),
  .ZN(_130_)
);

INV_X1 _220_ (
  .A(_130_),
  .ZN(_131_)
);

AOI21_X2 _221_ (
  .A(_098_),
  .B1(_128_),
  .B2(_131_),
  .ZN(_132_)
);

NAND2_X2 _222_ (
  .A1(_100_),
  .A2(_172_),
  .ZN(_133_)
);

INV_X1 _223_ (
  .A(_178_),
  .ZN(_134_)
);

NAND2_X4 _224_ (
  .A1(_134_),
  .A2(_104_),
  .ZN(_135_)
);

NAND3_X4 _225_ (
  .A1(_133_),
  .A2(_135_),
  .A3(_109_),
  .ZN(_136_)
);

NAND2_X4 _226_ (
  .A1(_100_),
  .A2(_103_),
  .ZN(_137_)
);

NAND2_X2 _227_ (
  .A1(_136_),
  .A2(_137_),
  .ZN(_138_)
);

INV_X1 _228_ (
  .A(y[1]),
  .ZN(_139_)
);

CLKBUF_X3 _229_ (
  .A(_139_),
  .Z(_140_)
);

NAND2_X1 _230_ (
  .A1(_138_),
  .A2(_140_),
  .ZN(_141_)
);

AOI21_X2 _231_ (
  .A(_122_),
  .B1(_132_),
  .B2(_141_),
  .ZN(_142_)
);

NAND2_X1 _232_ (
  .A1(_120_),
  .A2(_142_),
  .ZN(_143_)
);

NAND2_X1 _233_ (
  .A1(_122_),
  .A2(\coef[21] ),
  .ZN(_144_)
);

NAND2_X2 _234_ (
  .A1(_143_),
  .A2(_144_),
  .ZN(_000_)
);

NOR2_X1 _235_ (
  .A1(_121_),
  .A2(\coef[23] ),
  .ZN(_145_)
);

NAND2_X2 _236_ (
  .A1(_114_),
  .A2(_116_),
  .ZN(_146_)
);

NAND2_X4 _237_ (
  .A1(_146_),
  .A2(_127_),
  .ZN(_147_)
);

NAND3_X2 _238_ (
  .A1(_124_),
  .A2(_115_),
  .A3(_125_),
  .ZN(_148_)
);

NAND3_X1 _239_ (
  .A1(_147_),
  .A2(_148_),
  .A3(_140_),
  .ZN(_149_)
);

NAND2_X1 _240_ (
  .A1(_118_),
  .A2(_110_),
  .ZN(_150_)
);

AOI21_X1 _241_ (
  .A(_097_),
  .B1(_150_),
  .B2(_108_),
  .ZN(_151_)
);

AOI21_X1 _242_ (
  .A(_122_),
  .B1(_149_),
  .B2(_151_),
  .ZN(_152_)
);

NAND2_X2 _243_ (
  .A1(_137_),
  .A2(_129_),
  .ZN(_153_)
);

AOI21_X1 _244_ (
  .A(_098_),
  .B1(_153_),
  .B2(_140_),
  .ZN(_154_)
);

NAND2_X1 _245_ (
  .A1(_147_),
  .A2(_148_),
  .ZN(_155_)
);

OAI21_X1 _246_ (
  .A(_154_),
  .B1(_155_),
  .B2(_140_),
  .ZN(_156_)
);

AOI21_X2 _247_ (
  .A(_145_),
  .B1(_152_),
  .B2(_156_),
  .ZN(_001_)
);

NOR2_X1 _248_ (
  .A1(_121_),
  .A2(\coef[24] ),
  .ZN(_009_)
);

AOI21_X2 _249_ (
  .A(_107_),
  .B1(_166_),
  .B2(_127_),
  .ZN(_010_)
);

AOI21_X1 _250_ (
  .A(_097_),
  .B1(_148_),
  .B2(_010_),
  .ZN(_011_)
);

NAND2_X1 _251_ (
  .A1(_100_),
  .A2(_176_),
  .ZN(_012_)
);

NAND2_X4 _252_ (
  .A1(_101_),
  .A2(_104_),
  .ZN(_013_)
);

NAND3_X2 _253_ (
  .A1(_012_),
  .A2(_013_),
  .A3(_109_),
  .ZN(_014_)
);

NAND2_X1 _254_ (
  .A1(_167_),
  .A2(_127_),
  .ZN(_015_)
);

NAND3_X1 _255_ (
  .A1(_014_),
  .A2(_108_),
  .A3(_015_),
  .ZN(_016_)
);

AOI21_X1 _256_ (
  .A(_122_),
  .B1(_011_),
  .B2(_016_),
  .ZN(_017_)
);

NAND2_X1 _257_ (
  .A1(_147_),
  .A2(_131_),
  .ZN(_018_)
);

NAND2_X2 _258_ (
  .A1(_100_),
  .A2(_134_),
  .ZN(_019_)
);

NAND2_X4 _259_ (
  .A1(_104_),
  .A2(_172_),
  .ZN(_020_)
);

NAND3_X4 _260_ (
  .A1(_019_),
  .A2(_103_),
  .A3(_020_),
  .ZN(_021_)
);

AOI21_X2 _261_ (
  .A(_107_),
  .B1(_115_),
  .B2(x[1]),
  .ZN(_022_)
);

NAND2_X1 _262_ (
  .A1(_021_),
  .A2(_022_),
  .ZN(_023_)
);

NAND3_X1 _263_ (
  .A1(_018_),
  .A2(_023_),
  .A3(_097_),
  .ZN(_024_)
);

AOI21_X2 _264_ (
  .A(_009_),
  .B1(_017_),
  .B2(_024_),
  .ZN(_002_)
);

NAND3_X1 _265_ (
  .A1(_014_),
  .A2(_106_),
  .A3(_107_),
  .ZN(_025_)
);

NAND3_X1 _266_ (
  .A1(_124_),
  .A2(_103_),
  .A3(_125_),
  .ZN(_026_)
);

INV_X1 _267_ (
  .A(_170_),
  .ZN(_027_)
);

NAND2_X1 _268_ (
  .A1(_100_),
  .A2(_027_),
  .ZN(_028_)
);

NAND2_X4 _269_ (
  .A1(_104_),
  .A2(_180_),
  .ZN(_029_)
);

NAND3_X1 _270_ (
  .A1(_028_),
  .A2(_115_),
  .A3(_029_),
  .ZN(_030_)
);

NAND3_X1 _271_ (
  .A1(_026_),
  .A2(_030_),
  .A3(_139_),
  .ZN(_031_)
);

NAND2_X1 _272_ (
  .A1(_025_),
  .A2(_031_),
  .ZN(_032_)
);

NAND2_X1 _273_ (
  .A1(_032_),
  .A2(_097_),
  .ZN(_033_)
);

NAND2_X1 _274_ (
  .A1(_136_),
  .A2(_021_),
  .ZN(_034_)
);

NAND2_X1 _275_ (
  .A1(_034_),
  .A2(_140_),
  .ZN(_035_)
);

INV_X1 _276_ (
  .A(_168_),
  .ZN(_036_)
);

NAND2_X2 _277_ (
  .A1(_100_),
  .A2(_036_),
  .ZN(_037_)
);

NAND2_X4 _278_ (
  .A1(_104_),
  .A2(_182_),
  .ZN(_038_)
);

NAND3_X1 _279_ (
  .A1(_037_),
  .A2(_127_),
  .A3(_038_),
  .ZN(_039_)
);

NAND3_X1 _280_ (
  .A1(_117_),
  .A2(_039_),
  .A3(_108_),
  .ZN(_040_)
);

NAND3_X1 _281_ (
  .A1(_035_),
  .A2(_040_),
  .A3(_098_),
  .ZN(_041_)
);

NAND3_X1 _282_ (
  .A1(_033_),
  .A2(_041_),
  .A3(_121_),
  .ZN(_042_)
);

NAND2_X1 _283_ (
  .A1(_122_),
  .A2(\coef[10] ),
  .ZN(_043_)
);

NAND2_X1 _284_ (
  .A1(_042_),
  .A2(_043_),
  .ZN(_003_)
);

NOR2_X1 _285_ (
  .A1(_121_),
  .A2(\coef[26] ),
  .ZN(_044_)
);

AOI21_X1 _286_ (
  .A(_107_),
  .B1(_115_),
  .B2(_100_),
  .ZN(_045_)
);

AOI21_X2 _287_ (
  .A(_098_),
  .B1(_147_),
  .B2(_045_),
  .ZN(_046_)
);

NAND3_X1 _288_ (
  .A1(_133_),
  .A2(_135_),
  .A3(_127_),
  .ZN(_047_)
);

NAND3_X1 _289_ (
  .A1(_047_),
  .A2(_108_),
  .A3(_110_),
  .ZN(_048_)
);

AOI21_X2 _290_ (
  .A(_122_),
  .B1(_046_),
  .B2(_048_),
  .ZN(_049_)
);

NAND2_X1 _291_ (
  .A1(_104_),
  .A2(_127_),
  .ZN(_050_)
);

NAND3_X1 _292_ (
  .A1(_148_),
  .A2(_108_),
  .A3(_050_),
  .ZN(_051_)
);

NAND3_X1 _293_ (
  .A1(_102_),
  .A2(_115_),
  .A3(_105_),
  .ZN(_052_)
);

NAND3_X1 _294_ (
  .A1(_052_),
  .A2(_140_),
  .A3(_137_),
  .ZN(_053_)
);

NAND3_X1 _295_ (
  .A1(_051_),
  .A2(_053_),
  .A3(_098_),
  .ZN(_054_)
);

AOI21_X2 _296_ (
  .A(_044_),
  .B1(_049_),
  .B2(_054_),
  .ZN(_004_)
);

NAND2_X2 _297_ (
  .A1(_037_),
  .A2(_038_),
  .ZN(_055_)
);

NOR3_X2 _298_ (
  .A1(_055_),
  .A2(_103_),
  .A3(_107_),
  .ZN(_056_)
);

NAND2_X1 _299_ (
  .A1(_103_),
  .A2(x[1]),
  .ZN(_057_)
);

OAI21_X1 _300_ (
  .A(_097_),
  .B1(_057_),
  .B2(_107_),
  .ZN(_058_)
);

NOR2_X2 _301_ (
  .A1(_056_),
  .A2(_058_),
  .ZN(_059_)
);

XNOR2_X2 _302_ (
  .A(_099_),
  .B(_169_),
  .ZN(_060_)
);

INV_X2 _303_ (
  .A(_060_),
  .ZN(_061_)
);

NAND2_X2 _304_ (
  .A1(_061_),
  .A2(_115_),
  .ZN(_062_)
);

NAND3_X1 _305_ (
  .A1(_062_),
  .A2(_108_),
  .A3(_021_),
  .ZN(_063_)
);

NAND2_X2 _306_ (
  .A1(_059_),
  .A2(_063_),
  .ZN(_064_)
);

NAND2_X1 _307_ (
  .A1(_060_),
  .A2(_127_),
  .ZN(_065_)
);

NAND3_X1 _308_ (
  .A1(_065_),
  .A2(_140_),
  .A3(_014_),
  .ZN(_066_)
);

NAND3_X1 _309_ (
  .A1(_028_),
  .A2(_103_),
  .A3(_029_),
  .ZN(_067_)
);

OAI21_X1 _310_ (
  .A(_107_),
  .B1(_167_),
  .B2(_103_),
  .ZN(_068_)
);

INV_X1 _311_ (
  .A(_068_),
  .ZN(_069_)
);

AOI21_X1 _312_ (
  .A(_097_),
  .B1(_067_),
  .B2(_069_),
  .ZN(_070_)
);

NAND2_X1 _313_ (
  .A1(_066_),
  .A2(_070_),
  .ZN(_071_)
);

NAND2_X2 _314_ (
  .A1(_064_),
  .A2(_071_),
  .ZN(_072_)
);

NAND2_X2 _315_ (
  .A1(_072_),
  .A2(_121_),
  .ZN(_073_)
);

NAND2_X1 _316_ (
  .A1(_122_),
  .A2(\coef[13] ),
  .ZN(_074_)
);

NAND2_X2 _317_ (
  .A1(_073_),
  .A2(_074_),
  .ZN(_005_)
);

NOR2_X1 _318_ (
  .A1(_121_),
  .A2(\coef[28] ),
  .ZN(_075_)
);

NAND3_X1 _319_ (
  .A1(_062_),
  .A2(_108_),
  .A3(_057_),
  .ZN(_076_)
);

NAND2_X1 _320_ (
  .A1(_150_),
  .A2(_140_),
  .ZN(_077_)
);

NAND2_X1 _321_ (
  .A1(_076_),
  .A2(_077_),
  .ZN(_078_)
);

NAND2_X1 _322_ (
  .A1(_078_),
  .A2(_098_),
  .ZN(_079_)
);

NOR2_X1 _323_ (
  .A1(_153_),
  .A2(_140_),
  .ZN(_080_)
);

NOR2_X1 _324_ (
  .A1(_080_),
  .A2(_098_),
  .ZN(_081_)
);

OAI21_X1 _325_ (
  .A(_022_),
  .B1(_060_),
  .B2(_115_),
  .ZN(_082_)
);

AOI21_X2 _326_ (
  .A(_122_),
  .B1(_081_),
  .B2(_082_),
  .ZN(_083_)
);

AOI21_X2 _327_ (
  .A(_075_),
  .B1(_079_),
  .B2(_083_),
  .ZN(_006_)
);

NOR2_X1 _328_ (
  .A1(_121_),
  .A2(\coef[29] ),
  .ZN(_084_)
);

AOI21_X1 _329_ (
  .A(_098_),
  .B1(_065_),
  .B2(_131_),
  .ZN(_085_)
);

NAND3_X1 _330_ (
  .A1(_019_),
  .A2(_115_),
  .A3(_020_),
  .ZN(_086_)
);

NAND3_X1 _331_ (
  .A1(_106_),
  .A2(_086_),
  .A3(_140_),
  .ZN(_087_)
);

AOI21_X1 _332_ (
  .A(_122_),
  .B1(_085_),
  .B2(_087_),
  .ZN(_088_)
);

NAND3_X1 _333_ (
  .A1(_012_),
  .A2(_013_),
  .A3(_127_),
  .ZN(_089_)
);

NAND3_X1 _334_ (
  .A1(_136_),
  .A2(_089_),
  .A3(_108_),
  .ZN(_090_)
);

NAND2_X1 _335_ (
  .A1(_062_),
  .A2(_010_),
  .ZN(_091_)
);

NAND3_X1 _336_ (
  .A1(_090_),
  .A2(_098_),
  .A3(_091_),
  .ZN(_092_)
);

AOI21_X2 _337_ (
  .A(_084_),
  .B1(_088_),
  .B2(_092_),
  .ZN(_007_)
);

NOR2_X1 _338_ (
  .A1(_121_),
  .A2(\coef[30] ),
  .ZN(_093_)
);

OAI21_X2 _339_ (
  .A(_097_),
  .B1(_115_),
  .B2(_139_),
  .ZN(_094_)
);

OAI21_X1 _340_ (
  .A(_094_),
  .B1(_127_),
  .B2(_107_),
  .ZN(_095_)
);

XNOR2_X1 _341_ (
  .A(_095_),
  .B(_166_),
  .ZN(_096_)
);

AOI21_X2 _342_ (
  .A(_093_),
  .B1(_096_),
  .B2(_121_),
  .ZN(_008_)
);

HA_X1 _343_ (
  .A(_166_),
  .B(_167_),
  .CO(_168_),
  .S(_169_)
);

HA_X1 _344_ (
  .A(_166_),
  .B(_167_),
  .CO(_170_),
  .S(_171_)
);

HA_X1 _345_ (
  .A(_166_),
  .B(x[1]),
  .CO(_172_),
  .S(_173_)
);

HA_X1 _346_ (
  .A(_166_),
  .B(x[1]),
  .CO(_174_),
  .S(_175_)
);

HA_X1 _347_ (
  .A(x[0]),
  .B(_167_),
  .CO(_176_),
  .S(_177_)
);

HA_X1 _348_ (
  .A(x[0]),
  .B(_167_),
  .CO(_178_),
  .S(_179_)
);

HA_X1 _349_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_180_),
  .S(_181_)
);

HA_X1 _350_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_182_),
  .S(_183_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_165_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_164_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_163_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_162_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_161_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_160_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_159_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_158_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_157_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$ca051f171e86125a3bcf4bd090f5be774b98c04e\dctu

module \$paramod$cf6677181b8958913bf11288905dc7e6338a7bf5\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _110_ (
  .A(x[1]),
  .ZN(_033_)
);

NAND2_X1 _111_ (
  .A1(_033_),
  .A2(x[2]),
  .ZN(_034_)
);

INV_X2 _112_ (
  .A(x[2]),
  .ZN(_035_)
);

NAND2_X1 _113_ (
  .A1(_035_),
  .A2(x[1]),
  .ZN(_036_)
);

NAND2_X2 _114_ (
  .A1(_034_),
  .A2(_036_),
  .ZN(_037_)
);

BUF_X2 _115_ (
  .A(y[0]),
  .Z(_038_)
);

NAND2_X2 _116_ (
  .A1(_037_),
  .A2(_038_),
  .ZN(_039_)
);

NAND2_X2 _117_ (
  .A1(_035_),
  .A2(_033_),
  .ZN(_040_)
);

NAND2_X1 _118_ (
  .A1(x[2]),
  .A2(x[1]),
  .ZN(_041_)
);

NAND2_X4 _119_ (
  .A1(_040_),
  .A2(_041_),
  .ZN(_042_)
);

INV_X2 _120_ (
  .A(_038_),
  .ZN(_043_)
);

NAND2_X2 _121_ (
  .A1(_042_),
  .A2(_043_),
  .ZN(_044_)
);

BUF_X2 _122_ (
  .A(y[1]),
  .Z(_045_)
);

INV_X2 _123_ (
  .A(_045_),
  .ZN(_046_)
);

NAND3_X1 _124_ (
  .A1(_039_),
  .A2(_044_),
  .A3(_046_),
  .ZN(_047_)
);

INV_X1 _125_ (
  .A(x[0]),
  .ZN(_048_)
);

NAND2_X4 _126_ (
  .A1(_048_),
  .A2(_035_),
  .ZN(_049_)
);

NAND2_X2 _127_ (
  .A1(x[0]),
  .A2(x[2]),
  .ZN(_050_)
);

NAND2_X4 _128_ (
  .A1(_049_),
  .A2(_050_),
  .ZN(_051_)
);

NAND2_X2 _129_ (
  .A1(_051_),
  .A2(_043_),
  .ZN(_052_)
);

NAND3_X1 _130_ (
  .A1(_049_),
  .A2(_038_),
  .A3(_050_),
  .ZN(_053_)
);

NAND3_X1 _131_ (
  .A1(_052_),
  .A2(_053_),
  .A3(_045_),
  .ZN(_054_)
);

BUF_X1 _132_ (
  .A(y[2]),
  .Z(_055_)
);

BUF_X2 _133_ (
  .A(_055_),
  .Z(_056_)
);

NAND3_X1 _134_ (
  .A1(_047_),
  .A2(_054_),
  .A3(_056_),
  .ZN(_057_)
);

NAND3_X2 _135_ (
  .A1(_039_),
  .A2(_044_),
  .A3(_045_),
  .ZN(_058_)
);

NAND3_X1 _136_ (
  .A1(_052_),
  .A2(_053_),
  .A3(_046_),
  .ZN(_059_)
);

INV_X1 _137_ (
  .A(_056_),
  .ZN(_060_)
);

NAND3_X1 _138_ (
  .A1(_058_),
  .A2(_059_),
  .A3(_060_),
  .ZN(_061_)
);

BUF_X1 _139_ (
  .A(ena),
  .Z(_062_)
);

BUF_X1 _140_ (
  .A(_062_),
  .Z(_063_)
);

NAND3_X1 _141_ (
  .A1(_057_),
  .A2(_061_),
  .A3(_063_),
  .ZN(_064_)
);

INV_X1 _142_ (
  .A(_062_),
  .ZN(_065_)
);

NAND2_X1 _143_ (
  .A1(_065_),
  .A2(\coef[21] ),
  .ZN(_066_)
);

NAND2_X1 _144_ (
  .A1(_064_),
  .A2(_066_),
  .ZN(_000_)
);

NOR2_X1 _145_ (
  .A1(_062_),
  .A2(\coef[22] ),
  .ZN(_067_)
);

XNOR2_X1 _146_ (
  .A(_042_),
  .B(_056_),
  .ZN(_068_)
);

AOI21_X1 _147_ (
  .A(_067_),
  .B1(_068_),
  .B2(_063_),
  .ZN(_001_)
);

NAND2_X2 _148_ (
  .A1(_051_),
  .A2(_038_),
  .ZN(_069_)
);

NAND3_X1 _149_ (
  .A1(_040_),
  .A2(_043_),
  .A3(_041_),
  .ZN(_070_)
);

NAND2_X1 _150_ (
  .A1(_069_),
  .A2(_070_),
  .ZN(_071_)
);

NAND2_X1 _151_ (
  .A1(_071_),
  .A2(_046_),
  .ZN(_072_)
);

NAND3_X2 _152_ (
  .A1(_049_),
  .A2(_043_),
  .A3(_050_),
  .ZN(_073_)
);

NAND3_X1 _153_ (
  .A1(_069_),
  .A2(_073_),
  .A3(_045_),
  .ZN(_074_)
);

NAND3_X1 _154_ (
  .A1(_072_),
  .A2(_074_),
  .A3(_056_),
  .ZN(_075_)
);

NAND2_X1 _155_ (
  .A1(_042_),
  .A2(_038_),
  .ZN(_076_)
);

NAND2_X1 _156_ (
  .A1(_076_),
  .A2(_073_),
  .ZN(_077_)
);

NAND2_X1 _157_ (
  .A1(_077_),
  .A2(_045_),
  .ZN(_078_)
);

NAND3_X1 _158_ (
  .A1(_069_),
  .A2(_073_),
  .A3(_046_),
  .ZN(_079_)
);

NAND3_X1 _159_ (
  .A1(_078_),
  .A2(_079_),
  .A3(_060_),
  .ZN(_080_)
);

NAND3_X1 _160_ (
  .A1(_075_),
  .A2(_080_),
  .A3(_063_),
  .ZN(_081_)
);

NAND2_X1 _161_ (
  .A1(_065_),
  .A2(\coef[23] ),
  .ZN(_082_)
);

NAND2_X1 _162_ (
  .A1(_081_),
  .A2(_082_),
  .ZN(_002_)
);

AOI21_X1 _163_ (
  .A(_055_),
  .B1(_037_),
  .B2(_046_),
  .ZN(_083_)
);

AOI21_X1 _164_ (
  .A(_065_),
  .B1(_058_),
  .B2(_083_),
  .ZN(_084_)
);

NAND2_X2 _165_ (
  .A1(_042_),
  .A2(_045_),
  .ZN(_085_)
);

NAND3_X1 _166_ (
  .A1(_047_),
  .A2(_056_),
  .A3(_085_),
  .ZN(_086_)
);

NAND2_X1 _167_ (
  .A1(_084_),
  .A2(_086_),
  .ZN(_087_)
);

NAND2_X1 _168_ (
  .A1(_065_),
  .A2(\coef[24] ),
  .ZN(_088_)
);

NAND2_X1 _169_ (
  .A1(_087_),
  .A2(_088_),
  .ZN(_003_)
);

NAND3_X1 _170_ (
  .A1(_078_),
  .A2(_059_),
  .A3(_056_),
  .ZN(_089_)
);

NAND3_X1 _171_ (
  .A1(_072_),
  .A2(_054_),
  .A3(_060_),
  .ZN(_090_)
);

NAND3_X1 _172_ (
  .A1(_089_),
  .A2(_090_),
  .A3(_063_),
  .ZN(_091_)
);

NAND2_X1 _173_ (
  .A1(_065_),
  .A2(\coef[25] ),
  .ZN(_092_)
);

NAND2_X1 _174_ (
  .A1(_091_),
  .A2(_092_),
  .ZN(_004_)
);

NAND3_X1 _175_ (
  .A1(_039_),
  .A2(_073_),
  .A3(_046_),
  .ZN(_093_)
);

NAND3_X1 _176_ (
  .A1(_058_),
  .A2(_093_),
  .A3(_056_),
  .ZN(_094_)
);

NAND2_X1 _177_ (
  .A1(_051_),
  .A2(_045_),
  .ZN(_095_)
);

NAND2_X1 _178_ (
  .A1(_037_),
  .A2(_046_),
  .ZN(_096_)
);

NAND3_X1 _179_ (
  .A1(_095_),
  .A2(_096_),
  .A3(_038_),
  .ZN(_097_)
);

AOI21_X1 _180_ (
  .A(_055_),
  .B1(_037_),
  .B2(_043_),
  .ZN(_098_)
);

NAND2_X1 _181_ (
  .A1(_097_),
  .A2(_098_),
  .ZN(_099_)
);

NAND2_X1 _182_ (
  .A1(_094_),
  .A2(_099_),
  .ZN(_010_)
);

NAND2_X1 _183_ (
  .A1(_010_),
  .A2(_063_),
  .ZN(_011_)
);

NAND2_X1 _184_ (
  .A1(_065_),
  .A2(\coef[26] ),
  .ZN(_012_)
);

NAND2_X1 _185_ (
  .A1(_011_),
  .A2(_012_),
  .ZN(_005_)
);

OAI21_X1 _186_ (
  .A(_083_),
  .B1(_046_),
  .B2(_051_),
  .ZN(_013_)
);

NAND2_X1 _187_ (
  .A1(_051_),
  .A2(_046_),
  .ZN(_014_)
);

NAND2_X1 _188_ (
  .A1(_014_),
  .A2(_085_),
  .ZN(_015_)
);

INV_X2 _189_ (
  .A(_015_),
  .ZN(_016_)
);

NAND2_X1 _190_ (
  .A1(_016_),
  .A2(_056_),
  .ZN(_017_)
);

NAND3_X1 _191_ (
  .A1(_013_),
  .A2(_063_),
  .A3(_017_),
  .ZN(_018_)
);

INV_X1 _192_ (
  .A(\coef[27] ),
  .ZN(_019_)
);

OAI21_X1 _193_ (
  .A(_018_),
  .B1(_063_),
  .B2(_019_),
  .ZN(_006_)
);

NAND3_X1 _194_ (
  .A1(_054_),
  .A2(_079_),
  .A3(_056_),
  .ZN(_020_)
);

NAND3_X1 _195_ (
  .A1(_059_),
  .A2(_074_),
  .A3(_060_),
  .ZN(_021_)
);

NAND3_X1 _196_ (
  .A1(_020_),
  .A2(_021_),
  .A3(_063_),
  .ZN(_022_)
);

NAND2_X1 _197_ (
  .A1(_065_),
  .A2(\coef[28] ),
  .ZN(_023_)
);

NAND2_X1 _198_ (
  .A1(_022_),
  .A2(_023_),
  .ZN(_007_)
);

NAND2_X1 _199_ (
  .A1(_016_),
  .A2(_043_),
  .ZN(_024_)
);

AOI21_X1 _200_ (
  .A(_055_),
  .B1(_042_),
  .B2(_038_),
  .ZN(_025_)
);

AOI21_X2 _201_ (
  .A(_065_),
  .B1(_024_),
  .B2(_025_),
  .ZN(_026_)
);

NAND2_X1 _202_ (
  .A1(_071_),
  .A2(_045_),
  .ZN(_027_)
);

NAND3_X1 _203_ (
  .A1(_047_),
  .A2(_027_),
  .A3(_056_),
  .ZN(_028_)
);

NAND2_X1 _204_ (
  .A1(_026_),
  .A2(_028_),
  .ZN(_029_)
);

NAND2_X1 _205_ (
  .A1(_065_),
  .A2(\coef[15] ),
  .ZN(_030_)
);

NAND2_X1 _206_ (
  .A1(_029_),
  .A2(_030_),
  .ZN(_008_)
);

NAND3_X1 _207_ (
  .A1(_052_),
  .A2(_053_),
  .A3(_063_),
  .ZN(_031_)
);

INV_X1 _208_ (
  .A(\coef[30] ),
  .ZN(_032_)
);

OAI21_X1 _209_ (
  .A(_031_),
  .B1(_063_),
  .B2(_032_),
  .ZN(_009_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_109_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_108_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_107_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_106_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_105_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_104_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_103_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_102_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_101_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_100_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$cf6677181b8958913bf11288905dc7e6338a7bf5\dctu

module \$paramod$d348381a5c8d7c369f0c055d305d608d67b77e86\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _56_ (
  .A(y[0]),
  .ZN(_42_)
);

INV_X1 _57_ (
  .A(y[1]),
  .ZN(_43_)
);

BUF_X4 _58_ (
  .A(ena),
  .Z(_08_)
);

INV_X4 _59_ (
  .A(_08_),
  .ZN(_09_)
);

BUF_X16 _60_ (
  .A(_09_),
  .Z(_10_)
);

NAND2_X4 _61_ (
  .A1(_10_),
  .A2(\coef[21] ),
  .ZN(_11_)
);

BUF_X4 _62_ (
  .A(y[2]),
  .Z(_12_)
);

NAND2_X1 _63_ (
  .A1(_12_),
  .A2(_50_),
  .ZN(_13_)
);

NAND2_X1 _64_ (
  .A1(_13_),
  .A2(_08_),
  .ZN(_14_)
);

NOR2_X1 _65_ (
  .A1(_12_),
  .A2(_48_),
  .ZN(_15_)
);

OAI21_X2 _66_ (
  .A(_11_),
  .B1(_14_),
  .B2(_15_),
  .ZN(_00_)
);

NAND2_X4 _67_ (
  .A1(_10_),
  .A2(\coef[22] ),
  .ZN(_16_)
);

OAI21_X2 _68_ (
  .A(_16_),
  .B1(y[1]),
  .B2(_10_),
  .ZN(_01_)
);

NAND2_X4 _69_ (
  .A1(_10_),
  .A2(\coef[23] ),
  .ZN(_17_)
);

OAI21_X2 _70_ (
  .A(_17_),
  .B1(_12_),
  .B2(_10_),
  .ZN(_02_)
);

NAND2_X4 _71_ (
  .A1(_10_),
  .A2(\coef[14] ),
  .ZN(_18_)
);

OAI21_X2 _72_ (
  .A(_18_),
  .B1(_43_),
  .B2(_10_),
  .ZN(_03_)
);

NAND2_X4 _73_ (
  .A1(_10_),
  .A2(\coef[13] ),
  .ZN(_19_)
);

NAND2_X1 _74_ (
  .A1(_12_),
  .A2(_52_),
  .ZN(_20_)
);

NAND2_X1 _75_ (
  .A1(_20_),
  .A2(_08_),
  .ZN(_21_)
);

NOR2_X1 _76_ (
  .A1(_12_),
  .A2(_46_),
  .ZN(_22_)
);

OAI21_X2 _77_ (
  .A(_19_),
  .B1(_21_),
  .B2(_22_),
  .ZN(_04_)
);

NAND2_X1 _78_ (
  .A1(_09_),
  .A2(\coef[28] ),
  .ZN(_23_)
);

NAND2_X1 _79_ (
  .A1(_12_),
  .A2(_44_),
  .ZN(_24_)
);

NAND2_X1 _80_ (
  .A1(_24_),
  .A2(_08_),
  .ZN(_25_)
);

NOR2_X1 _81_ (
  .A1(_12_),
  .A2(_54_),
  .ZN(_26_)
);

OAI21_X1 _82_ (
  .A(_23_),
  .B1(_25_),
  .B2(_26_),
  .ZN(_05_)
);

INV_X1 _83_ (
  .A(_12_),
  .ZN(_27_)
);

INV_X1 _84_ (
  .A(_45_),
  .ZN(_28_)
);

NAND2_X1 _85_ (
  .A1(_27_),
  .A2(_28_),
  .ZN(_29_)
);

NAND2_X1 _86_ (
  .A1(_12_),
  .A2(_45_),
  .ZN(_30_)
);

NAND3_X1 _87_ (
  .A1(_29_),
  .A2(_08_),
  .A3(_30_),
  .ZN(_31_)
);

NAND2_X4 _88_ (
  .A1(_10_),
  .A2(\coef[15] ),
  .ZN(_32_)
);

NAND2_X2 _89_ (
  .A1(_31_),
  .A2(_32_),
  .ZN(_06_)
);

NAND2_X1 _90_ (
  .A1(_09_),
  .A2(\coef[12] ),
  .ZN(_33_)
);

OAI21_X2 _91_ (
  .A(_33_),
  .B1(_42_),
  .B2(_10_),
  .ZN(_07_)
);

HA_X1 _92_ (
  .A(_42_),
  .B(_43_),
  .CO(_44_),
  .S(_45_)
);

HA_X1 _93_ (
  .A(_42_),
  .B(_43_),
  .CO(_46_),
  .S(_47_)
);

HA_X1 _94_ (
  .A(_42_),
  .B(y[1]),
  .CO(_48_),
  .S(_49_)
);

HA_X1 _95_ (
  .A(y[0]),
  .B(_43_),
  .CO(_50_),
  .S(_51_)
);

HA_X1 _96_ (
  .A(y[0]),
  .B(y[1]),
  .CO(_52_),
  .S(_53_)
);

HA_X1 _97_ (
  .A(y[0]),
  .B(y[1]),
  .CO(_54_),
  .S(_55_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_41_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_01_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_40_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_02_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_39_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_03_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_38_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_04_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_37_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_05_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_36_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_06_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_35_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_07_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_34_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$d348381a5c8d7c369f0c055d305d608d67b77e86\dctu

module \$paramod$da3415da01ee30cd3fa431ef7b8104a7c6ed9a24\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _174_ (
  .A(x[1]),
  .ZN(_157_)
);

INV_X1 _175_ (
  .A(x[0]),
  .ZN(_156_)
);

BUF_X1 _176_ (
  .A(ena),
  .Z(_090_)
);

NOR2_X1 _177_ (
  .A1(\coef[21] ),
  .A2(_090_),
  .ZN(_091_)
);

BUF_X8 _178_ (
  .A(y[0]),
  .Z(_092_)
);

INV_X8 _179_ (
  .A(_092_),
  .ZN(_093_)
);

BUF_X8 _180_ (
  .A(x[2]),
  .Z(_094_)
);

NOR2_X4 _181_ (
  .A1(_093_),
  .A2(_094_),
  .ZN(_095_)
);

INV_X2 _182_ (
  .A(_095_),
  .ZN(_096_)
);

NAND2_X2 _183_ (
  .A1(_093_),
  .A2(x[1]),
  .ZN(_097_)
);

NAND2_X2 _184_ (
  .A1(_096_),
  .A2(_097_),
  .ZN(_098_)
);

BUF_X4 _185_ (
  .A(y[1]),
  .Z(_099_)
);

INV_X1 _186_ (
  .A(_099_),
  .ZN(_100_)
);

NAND2_X2 _187_ (
  .A1(_098_),
  .A2(_100_),
  .ZN(_101_)
);

NOR2_X2 _188_ (
  .A1(_094_),
  .A2(_092_),
  .ZN(_102_)
);

INV_X1 _189_ (
  .A(_102_),
  .ZN(_103_)
);

NAND2_X1 _190_ (
  .A1(_092_),
  .A2(x[1]),
  .ZN(_104_)
);

NAND3_X1 _191_ (
  .A1(_103_),
  .A2(_099_),
  .A3(_104_),
  .ZN(_105_)
);

NAND2_X2 _192_ (
  .A1(_101_),
  .A2(_105_),
  .ZN(_106_)
);

BUF_X4 _193_ (
  .A(y[2]),
  .Z(_107_)
);

INV_X4 _194_ (
  .A(_107_),
  .ZN(_108_)
);

XNOR2_X2 _195_ (
  .A(_106_),
  .B(_108_),
  .ZN(_109_)
);

BUF_X2 _196_ (
  .A(_090_),
  .Z(_110_)
);

AOI21_X2 _197_ (
  .A(_091_),
  .B1(_109_),
  .B2(_110_),
  .ZN(_000_)
);

NOR2_X1 _198_ (
  .A1(_110_),
  .A2(\coef[22] ),
  .ZN(_111_)
);

NAND2_X1 _199_ (
  .A1(_092_),
  .A2(_107_),
  .ZN(_112_)
);

INV_X1 _200_ (
  .A(_112_),
  .ZN(_113_)
);

NOR2_X1 _201_ (
  .A1(_092_),
  .A2(_107_),
  .ZN(_114_)
);

NOR2_X2 _202_ (
  .A1(_113_),
  .A2(_114_),
  .ZN(_115_)
);

XNOR2_X1 _203_ (
  .A(_115_),
  .B(_156_),
  .ZN(_116_)
);

AOI21_X1 _204_ (
  .A(_111_),
  .B1(_116_),
  .B2(_110_),
  .ZN(_001_)
);

NOR2_X1 _205_ (
  .A1(_110_),
  .A2(\coef[23] ),
  .ZN(_117_)
);

INV_X1 _206_ (
  .A(_090_),
  .ZN(_118_)
);

BUF_X8 _207_ (
  .A(_092_),
  .Z(_119_)
);

AOI21_X2 _208_ (
  .A(_099_),
  .B1(_157_),
  .B2(_119_),
  .ZN(_120_)
);

BUF_X16 _209_ (
  .A(_094_),
  .Z(_121_)
);

NAND2_X2 _210_ (
  .A1(_121_),
  .A2(_162_),
  .ZN(_122_)
);

OAI21_X2 _211_ (
  .A(_122_),
  .B1(_121_),
  .B2(_168_),
  .ZN(_123_)
);

OAI21_X1 _212_ (
  .A(_120_),
  .B1(_123_),
  .B2(_119_),
  .ZN(_124_)
);

NAND2_X2 _213_ (
  .A1(_121_),
  .A2(_164_),
  .ZN(_125_)
);

OAI21_X1 _214_ (
  .A(_125_),
  .B1(_121_),
  .B2(_166_),
  .ZN(_126_)
);

NAND2_X1 _215_ (
  .A1(_126_),
  .A2(_113_),
  .ZN(_127_)
);

NAND2_X1 _216_ (
  .A1(_097_),
  .A2(_099_),
  .ZN(_128_)
);

NAND2_X1 _217_ (
  .A1(_128_),
  .A2(_107_),
  .ZN(_129_)
);

NAND2_X1 _218_ (
  .A1(_127_),
  .A2(_129_),
  .ZN(_130_)
);

AOI21_X1 _219_ (
  .A(_118_),
  .B1(_124_),
  .B2(_130_),
  .ZN(_131_)
);

OAI21_X1 _220_ (
  .A(_120_),
  .B1(_126_),
  .B2(_119_),
  .ZN(_132_)
);

NAND2_X1 _221_ (
  .A1(_123_),
  .A2(_119_),
  .ZN(_133_)
);

INV_X1 _222_ (
  .A(_128_),
  .ZN(_134_)
);

NAND2_X1 _223_ (
  .A1(_133_),
  .A2(_134_),
  .ZN(_135_)
);

NAND2_X1 _224_ (
  .A1(_132_),
  .A2(_135_),
  .ZN(_136_)
);

NAND2_X1 _225_ (
  .A1(_136_),
  .A2(_108_),
  .ZN(_137_)
);

AOI21_X2 _226_ (
  .A(_117_),
  .B1(_131_),
  .B2(_137_),
  .ZN(_002_)
);

NAND2_X1 _227_ (
  .A1(_121_),
  .A2(_168_),
  .ZN(_138_)
);

OAI21_X1 _228_ (
  .A(_138_),
  .B1(_121_),
  .B2(_162_),
  .ZN(_139_)
);

OR2_X1 _229_ (
  .A1(_139_),
  .A2(_115_),
  .ZN(_140_)
);

INV_X4 _230_ (
  .A(_094_),
  .ZN(_141_)
);

NAND2_X1 _231_ (
  .A1(_141_),
  .A2(_164_),
  .ZN(_142_)
);

OR2_X1 _232_ (
  .A1(_141_),
  .A2(_166_),
  .ZN(_143_)
);

NAND3_X1 _233_ (
  .A1(_115_),
  .A2(_142_),
  .A3(_143_),
  .ZN(_144_)
);

NAND3_X1 _234_ (
  .A1(_140_),
  .A2(_144_),
  .A3(_110_),
  .ZN(_145_)
);

INV_X1 _235_ (
  .A(\coef[24] ),
  .ZN(_010_)
);

OAI21_X1 _236_ (
  .A(_145_),
  .B1(_110_),
  .B2(_010_),
  .ZN(_003_)
);

NOR2_X1 _237_ (
  .A1(_110_),
  .A2(\coef[25] ),
  .ZN(_011_)
);

NAND2_X2 _238_ (
  .A1(_141_),
  .A2(_170_),
  .ZN(_012_)
);

INV_X1 _239_ (
  .A(_160_),
  .ZN(_013_)
);

NAND2_X1 _240_ (
  .A1(_013_),
  .A2(_094_),
  .ZN(_014_)
);

NAND3_X1 _241_ (
  .A1(_012_),
  .A2(_014_),
  .A3(_119_),
  .ZN(_015_)
);

NAND2_X1 _242_ (
  .A1(_015_),
  .A2(_103_),
  .ZN(_016_)
);

NAND2_X1 _243_ (
  .A1(_108_),
  .A2(_099_),
  .ZN(_017_)
);

INV_X1 _244_ (
  .A(_017_),
  .ZN(_018_)
);

NAND2_X1 _245_ (
  .A1(_016_),
  .A2(_018_),
  .ZN(_019_)
);

INV_X1 _246_ (
  .A(_172_),
  .ZN(_020_)
);

NAND2_X2 _247_ (
  .A1(_141_),
  .A2(_020_),
  .ZN(_021_)
);

NAND2_X1 _248_ (
  .A1(_094_),
  .A2(_158_),
  .ZN(_022_)
);

NAND3_X1 _249_ (
  .A1(_021_),
  .A2(_119_),
  .A3(_022_),
  .ZN(_023_)
);

NAND2_X1 _250_ (
  .A1(_093_),
  .A2(_121_),
  .ZN(_024_)
);

NAND2_X1 _251_ (
  .A1(_023_),
  .A2(_024_),
  .ZN(_025_)
);

NAND2_X1 _252_ (
  .A1(_099_),
  .A2(_107_),
  .ZN(_026_)
);

INV_X1 _253_ (
  .A(_026_),
  .ZN(_027_)
);

NAND2_X1 _254_ (
  .A1(_025_),
  .A2(_027_),
  .ZN(_028_)
);

NAND2_X1 _255_ (
  .A1(_019_),
  .A2(_028_),
  .ZN(_029_)
);

NOR2_X2 _256_ (
  .A1(_108_),
  .A2(y[1]),
  .ZN(_030_)
);

INV_X1 _257_ (
  .A(_030_),
  .ZN(_031_)
);

NAND3_X1 _258_ (
  .A1(_012_),
  .A2(_014_),
  .A3(_093_),
  .ZN(_032_)
);

AOI21_X1 _259_ (
  .A(_031_),
  .B1(_032_),
  .B2(_096_),
  .ZN(_033_)
);

NOR2_X1 _260_ (
  .A1(_029_),
  .A2(_033_),
  .ZN(_034_)
);

NAND3_X1 _261_ (
  .A1(_021_),
  .A2(_093_),
  .A3(_022_),
  .ZN(_035_)
);

NAND2_X1 _262_ (
  .A1(_094_),
  .A2(_092_),
  .ZN(_036_)
);

NAND2_X1 _263_ (
  .A1(_035_),
  .A2(_036_),
  .ZN(_037_)
);

NOR2_X1 _264_ (
  .A1(_099_),
  .A2(_107_),
  .ZN(_038_)
);

AOI21_X1 _265_ (
  .A(_118_),
  .B1(_037_),
  .B2(_038_),
  .ZN(_039_)
);

AOI21_X2 _266_ (
  .A(_011_),
  .B1(_034_),
  .B2(_039_),
  .ZN(_004_)
);

NAND2_X1 _267_ (
  .A1(_118_),
  .A2(\coef[26] ),
  .ZN(_040_)
);

NAND2_X1 _268_ (
  .A1(_141_),
  .A2(_013_),
  .ZN(_041_)
);

NAND2_X1 _269_ (
  .A1(_121_),
  .A2(_170_),
  .ZN(_042_)
);

NAND2_X1 _270_ (
  .A1(_041_),
  .A2(_042_),
  .ZN(_043_)
);

NAND2_X1 _271_ (
  .A1(_043_),
  .A2(_093_),
  .ZN(_044_)
);

NAND2_X1 _272_ (
  .A1(_036_),
  .A2(_099_),
  .ZN(_045_)
);

INV_X1 _273_ (
  .A(_045_),
  .ZN(_046_)
);

NAND2_X1 _274_ (
  .A1(_044_),
  .A2(_046_),
  .ZN(_047_)
);

NAND2_X1 _275_ (
  .A1(_141_),
  .A2(_158_),
  .ZN(_048_)
);

NAND2_X2 _276_ (
  .A1(_020_),
  .A2(_121_),
  .ZN(_049_)
);

NAND2_X2 _277_ (
  .A1(_048_),
  .A2(_049_),
  .ZN(_050_)
);

NAND2_X1 _278_ (
  .A1(_050_),
  .A2(_119_),
  .ZN(_051_)
);

NOR2_X1 _279_ (
  .A1(_102_),
  .A2(_099_),
  .ZN(_052_)
);

NAND2_X1 _280_ (
  .A1(_051_),
  .A2(_052_),
  .ZN(_053_)
);

NAND3_X1 _281_ (
  .A1(_047_),
  .A2(_053_),
  .A3(_108_),
  .ZN(_054_)
);

NAND2_X1 _282_ (
  .A1(_054_),
  .A2(_110_),
  .ZN(_055_)
);

OAI21_X1 _283_ (
  .A(_052_),
  .B1(_043_),
  .B2(_093_),
  .ZN(_056_)
);

OAI21_X1 _284_ (
  .A(_046_),
  .B1(_050_),
  .B2(_119_),
  .ZN(_057_)
);

AOI21_X1 _285_ (
  .A(_108_),
  .B1(_056_),
  .B2(_057_),
  .ZN(_058_)
);

OAI21_X2 _286_ (
  .A(_040_),
  .B1(_055_),
  .B2(_058_),
  .ZN(_005_)
);

OR2_X4 _287_ (
  .A1(_159_),
  .A2(_094_),
  .ZN(_059_)
);

NAND2_X1 _288_ (
  .A1(_094_),
  .A2(_159_),
  .ZN(_060_)
);

NAND2_X2 _289_ (
  .A1(_059_),
  .A2(_060_),
  .ZN(_061_)
);

NAND2_X2 _290_ (
  .A1(_061_),
  .A2(_093_),
  .ZN(_062_)
);

AOI21_X1 _291_ (
  .A(_099_),
  .B1(_156_),
  .B2(_119_),
  .ZN(_063_)
);

NAND2_X2 _292_ (
  .A1(_062_),
  .A2(_063_),
  .ZN(_064_)
);

NAND3_X1 _293_ (
  .A1(_059_),
  .A2(_119_),
  .A3(_060_),
  .ZN(_065_)
);

OAI21_X1 _294_ (
  .A(y[1]),
  .B1(_156_),
  .B2(_092_),
  .ZN(_066_)
);

INV_X1 _295_ (
  .A(_066_),
  .ZN(_067_)
);

NAND2_X1 _296_ (
  .A1(_065_),
  .A2(_067_),
  .ZN(_068_)
);

NAND2_X1 _297_ (
  .A1(_064_),
  .A2(_068_),
  .ZN(_069_)
);

NAND2_X1 _298_ (
  .A1(_069_),
  .A2(_108_),
  .ZN(_070_)
);

NAND3_X1 _299_ (
  .A1(_064_),
  .A2(_068_),
  .A3(_107_),
  .ZN(_071_)
);

NAND3_X1 _300_ (
  .A1(_070_),
  .A2(_071_),
  .A3(_110_),
  .ZN(_072_)
);

NAND2_X1 _301_ (
  .A1(_118_),
  .A2(\coef[27] ),
  .ZN(_073_)
);

NAND2_X1 _302_ (
  .A1(_072_),
  .A2(_073_),
  .ZN(_006_)
);

NOR2_X1 _303_ (
  .A1(_090_),
  .A2(\coef[28] ),
  .ZN(_074_)
);

NAND2_X2 _304_ (
  .A1(_031_),
  .A2(_017_),
  .ZN(_075_)
);

XNOR2_X1 _305_ (
  .A(_075_),
  .B(_157_),
  .ZN(_076_)
);

AOI21_X1 _306_ (
  .A(_074_),
  .B1(_076_),
  .B2(_110_),
  .ZN(_007_)
);

NOR2_X1 _307_ (
  .A1(_090_),
  .A2(\coef[15] ),
  .ZN(_077_)
);

NAND2_X1 _308_ (
  .A1(_035_),
  .A2(_096_),
  .ZN(_078_)
);

NAND2_X1 _309_ (
  .A1(_078_),
  .A2(_030_),
  .ZN(_079_)
);

NAND2_X1 _310_ (
  .A1(_023_),
  .A2(_103_),
  .ZN(_080_)
);

NAND2_X1 _311_ (
  .A1(_080_),
  .A2(_018_),
  .ZN(_081_)
);

NAND2_X1 _312_ (
  .A1(_079_),
  .A2(_081_),
  .ZN(_082_)
);

INV_X1 _313_ (
  .A(_038_),
  .ZN(_083_)
);

AOI21_X1 _314_ (
  .A(_083_),
  .B1(_032_),
  .B2(_036_),
  .ZN(_084_)
);

NOR2_X2 _315_ (
  .A1(_082_),
  .A2(_084_),
  .ZN(_085_)
);

NAND2_X1 _316_ (
  .A1(_015_),
  .A2(_024_),
  .ZN(_086_)
);

AOI21_X1 _317_ (
  .A(_118_),
  .B1(_086_),
  .B2(_027_),
  .ZN(_087_)
);

AOI21_X2 _318_ (
  .A(_077_),
  .B1(_085_),
  .B2(_087_),
  .ZN(_008_)
);

NAND2_X1 _319_ (
  .A1(_118_),
  .A2(\coef[30] ),
  .ZN(_088_)
);

XNOR2_X1 _320_ (
  .A(_075_),
  .B(_121_),
  .ZN(_089_)
);

OAI21_X1 _321_ (
  .A(_088_),
  .B1(_089_),
  .B2(_118_),
  .ZN(_009_)
);

HA_X1 _322_ (
  .A(_156_),
  .B(_157_),
  .CO(_158_),
  .S(_159_)
);

HA_X1 _323_ (
  .A(_156_),
  .B(_157_),
  .CO(_160_),
  .S(_161_)
);

HA_X1 _324_ (
  .A(_156_),
  .B(x[1]),
  .CO(_162_),
  .S(_163_)
);

HA_X1 _325_ (
  .A(_156_),
  .B(x[1]),
  .CO(_164_),
  .S(_165_)
);

HA_X1 _326_ (
  .A(x[0]),
  .B(_157_),
  .CO(_166_),
  .S(_167_)
);

HA_X1 _327_ (
  .A(x[0]),
  .B(_157_),
  .CO(_168_),
  .S(_169_)
);

HA_X1 _328_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_170_),
  .S(_171_)
);

HA_X1 _329_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_172_),
  .S(_173_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_155_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_154_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_153_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_152_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_151_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_150_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_149_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_148_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_147_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_146_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$da3415da01ee30cd3fa431ef7b8104a7c6ed9a24\dctu

module \$paramod$e2471d3acfddfd8f107137e4952b02d9e7720f44\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[21] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[26] ;
wire \coef[28] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _189_ (
  .A(x[1]),
  .ZN(_172_)
);

INV_X1 _190_ (
  .A(x[0]),
  .ZN(_171_)
);

BUF_X2 _191_ (
  .A(ena),
  .Z(_102_)
);

INV_X1 _192_ (
  .A(_102_),
  .ZN(_103_)
);

NAND2_X1 _193_ (
  .A1(_103_),
  .A2(\coef[21] ),
  .ZN(_104_)
);

BUF_X4 _194_ (
  .A(x[2]),
  .Z(_105_)
);

INV_X4 _195_ (
  .A(_105_),
  .ZN(_106_)
);

INV_X1 _196_ (
  .A(_173_),
  .ZN(_107_)
);

NAND2_X1 _197_ (
  .A1(_106_),
  .A2(_107_),
  .ZN(_108_)
);

BUF_X4 _198_ (
  .A(y[0]),
  .Z(_109_)
);

INV_X8 _199_ (
  .A(_109_),
  .ZN(_110_)
);

NAND2_X1 _200_ (
  .A1(_105_),
  .A2(_187_),
  .ZN(_111_)
);

NAND3_X2 _201_ (
  .A1(_108_),
  .A2(_110_),
  .A3(_111_),
  .ZN(_112_)
);

BUF_X2 _202_ (
  .A(y[1]),
  .Z(_113_)
);

INV_X1 _203_ (
  .A(_113_),
  .ZN(_114_)
);

NAND2_X1 _204_ (
  .A1(_172_),
  .A2(_109_),
  .ZN(_115_)
);

NAND3_X1 _205_ (
  .A1(_112_),
  .A2(_114_),
  .A3(_115_),
  .ZN(_116_)
);

INV_X1 _206_ (
  .A(_174_),
  .ZN(_117_)
);

NAND2_X1 _207_ (
  .A1(_117_),
  .A2(_105_),
  .ZN(_118_)
);

NAND2_X4 _208_ (
  .A1(_106_),
  .A2(_174_),
  .ZN(_119_)
);

NAND2_X2 _209_ (
  .A1(_118_),
  .A2(_119_),
  .ZN(_120_)
);

BUF_X16 _210_ (
  .A(_110_),
  .Z(_121_)
);

NAND3_X1 _211_ (
  .A1(_120_),
  .A2(_121_),
  .A3(_113_),
  .ZN(_122_)
);

NAND2_X1 _212_ (
  .A1(_116_),
  .A2(_122_),
  .ZN(_123_)
);

NAND2_X1 _213_ (
  .A1(_106_),
  .A2(_181_),
  .ZN(_124_)
);

INV_X1 _214_ (
  .A(_179_),
  .ZN(_125_)
);

BUF_X8 _215_ (
  .A(_105_),
  .Z(_126_)
);

NAND2_X2 _216_ (
  .A1(_125_),
  .A2(_126_),
  .ZN(_127_)
);

AND2_X2 _217_ (
  .A1(_124_),
  .A2(_127_),
  .ZN(_128_)
);

BUF_X4 _218_ (
  .A(_109_),
  .Z(_129_)
);

BUF_X2 _219_ (
  .A(_113_),
  .Z(_130_)
);

NAND3_X1 _220_ (
  .A1(_128_),
  .A2(_129_),
  .A3(_130_),
  .ZN(_131_)
);

BUF_X2 _221_ (
  .A(y[2]),
  .Z(_132_)
);

INV_X1 _222_ (
  .A(_132_),
  .ZN(_133_)
);

BUF_X2 _223_ (
  .A(_133_),
  .Z(_134_)
);

NAND2_X1 _224_ (
  .A1(_131_),
  .A2(_134_),
  .ZN(_135_)
);

OAI21_X1 _225_ (
  .A(_102_),
  .B1(_123_),
  .B2(_135_),
  .ZN(_136_)
);

INV_X1 _226_ (
  .A(_175_),
  .ZN(_137_)
);

NAND2_X1 _227_ (
  .A1(_106_),
  .A2(_137_),
  .ZN(_138_)
);

NAND2_X2 _228_ (
  .A1(_126_),
  .A2(_185_),
  .ZN(_139_)
);

NAND2_X2 _229_ (
  .A1(_138_),
  .A2(_139_),
  .ZN(_140_)
);

NAND2_X2 _230_ (
  .A1(_140_),
  .A2(_129_),
  .ZN(_141_)
);

NAND2_X2 _231_ (
  .A1(_110_),
  .A2(x[1]),
  .ZN(_142_)
);

NAND2_X1 _232_ (
  .A1(_142_),
  .A2(_113_),
  .ZN(_143_)
);

INV_X1 _233_ (
  .A(_143_),
  .ZN(_144_)
);

AOI21_X1 _234_ (
  .A(_134_),
  .B1(_141_),
  .B2(_144_),
  .ZN(_145_)
);

INV_X1 _235_ (
  .A(_183_),
  .ZN(_146_)
);

NAND2_X2 _236_ (
  .A1(_106_),
  .A2(_146_),
  .ZN(_147_)
);

NAND2_X4 _237_ (
  .A1(_126_),
  .A2(_177_),
  .ZN(_148_)
);

NAND2_X1 _238_ (
  .A1(_147_),
  .A2(_148_),
  .ZN(_149_)
);

NAND2_X1 _239_ (
  .A1(_149_),
  .A2(_121_),
  .ZN(_150_)
);

NAND2_X2 _240_ (
  .A1(_120_),
  .A2(_129_),
  .ZN(_151_)
);

NAND3_X1 _241_ (
  .A1(_150_),
  .A2(_151_),
  .A3(_114_),
  .ZN(_152_)
);

AND2_X1 _242_ (
  .A1(_145_),
  .A2(_152_),
  .ZN(_153_)
);

OAI21_X2 _243_ (
  .A(_104_),
  .B1(_136_),
  .B2(_153_),
  .ZN(_000_)
);

NAND2_X1 _244_ (
  .A1(_109_),
  .A2(_113_),
  .ZN(_154_)
);

AOI21_X1 _245_ (
  .A(_154_),
  .B1(_108_),
  .B2(_111_),
  .ZN(_155_)
);

INV_X1 _246_ (
  .A(_142_),
  .ZN(_156_)
);

NOR3_X1 _247_ (
  .A1(_155_),
  .A2(_134_),
  .A3(_156_),
  .ZN(_157_)
);

NAND3_X4 _248_ (
  .A1(_147_),
  .A2(_109_),
  .A3(_148_),
  .ZN(_158_)
);

OR2_X4 _249_ (
  .A1(_158_),
  .A2(_130_),
  .ZN(_159_)
);

AOI21_X2 _250_ (
  .A(_103_),
  .B1(_157_),
  .B2(_159_),
  .ZN(_160_)
);

OAI21_X1 _251_ (
  .A(_115_),
  .B1(_140_),
  .B2(_129_),
  .ZN(_161_)
);

NAND2_X1 _252_ (
  .A1(_161_),
  .A2(_114_),
  .ZN(_009_)
);

NAND3_X2 _253_ (
  .A1(_124_),
  .A2(_127_),
  .A3(_110_),
  .ZN(_010_)
);

NAND2_X1 _254_ (
  .A1(_010_),
  .A2(_115_),
  .ZN(_011_)
);

NAND2_X1 _255_ (
  .A1(_011_),
  .A2(_130_),
  .ZN(_012_)
);

NAND3_X1 _256_ (
  .A1(_009_),
  .A2(_012_),
  .A3(_134_),
  .ZN(_013_)
);

NAND2_X1 _257_ (
  .A1(_160_),
  .A2(_013_),
  .ZN(_014_)
);

NAND2_X1 _258_ (
  .A1(_103_),
  .A2(\coef[23] ),
  .ZN(_015_)
);

NAND2_X1 _259_ (
  .A1(_014_),
  .A2(_015_),
  .ZN(_001_)
);

NOR2_X1 _260_ (
  .A1(_102_),
  .A2(\coef[24] ),
  .ZN(_016_)
);

NAND2_X1 _261_ (
  .A1(_106_),
  .A2(_177_),
  .ZN(_017_)
);

NAND2_X1 _262_ (
  .A1(_146_),
  .A2(_126_),
  .ZN(_018_)
);

NAND3_X1 _263_ (
  .A1(_017_),
  .A2(_018_),
  .A3(_121_),
  .ZN(_019_)
);

NAND3_X1 _264_ (
  .A1(_019_),
  .A2(_158_),
  .A3(_113_),
  .ZN(_020_)
);

AOI21_X1 _265_ (
  .A(_113_),
  .B1(_121_),
  .B2(_126_),
  .ZN(_021_)
);

AOI21_X1 _266_ (
  .A(_132_),
  .B1(_021_),
  .B2(_115_),
  .ZN(_022_)
);

AOI21_X1 _267_ (
  .A(_103_),
  .B1(_020_),
  .B2(_022_),
  .ZN(_023_)
);

NAND2_X1 _268_ (
  .A1(_106_),
  .A2(_125_),
  .ZN(_024_)
);

NAND2_X1 _269_ (
  .A1(_126_),
  .A2(_181_),
  .ZN(_025_)
);

NAND3_X1 _270_ (
  .A1(_024_),
  .A2(_109_),
  .A3(_025_),
  .ZN(_026_)
);

NAND3_X1 _271_ (
  .A1(_010_),
  .A2(_026_),
  .A3(_114_),
  .ZN(_027_)
);

NOR2_X2 _272_ (
  .A1(_110_),
  .A2(_126_),
  .ZN(_028_)
);

INV_X1 _273_ (
  .A(_028_),
  .ZN(_029_)
);

NAND3_X1 _274_ (
  .A1(_029_),
  .A2(_130_),
  .A3(_142_),
  .ZN(_030_)
);

NAND3_X1 _275_ (
  .A1(_027_),
  .A2(_132_),
  .A3(_030_),
  .ZN(_031_)
);

AOI21_X1 _276_ (
  .A(_016_),
  .B1(_023_),
  .B2(_031_),
  .ZN(_002_)
);

NOR2_X1 _277_ (
  .A1(_102_),
  .A2(\coef[10] ),
  .ZN(_032_)
);

INV_X1 _278_ (
  .A(_154_),
  .ZN(_033_)
);

AOI21_X1 _279_ (
  .A(_133_),
  .B1(_033_),
  .B2(_172_),
  .ZN(_034_)
);

NAND2_X1 _280_ (
  .A1(_122_),
  .A2(_034_),
  .ZN(_035_)
);

INV_X1 _281_ (
  .A(_035_),
  .ZN(_036_)
);

NAND2_X1 _282_ (
  .A1(_129_),
  .A2(x[0]),
  .ZN(_037_)
);

NAND2_X1 _283_ (
  .A1(_021_),
  .A2(_037_),
  .ZN(_038_)
);

AOI21_X1 _284_ (
  .A(_103_),
  .B1(_036_),
  .B2(_038_),
  .ZN(_039_)
);

AOI21_X1 _285_ (
  .A(_113_),
  .B1(_172_),
  .B2(_121_),
  .ZN(_040_)
);

AOI21_X2 _286_ (
  .A(_132_),
  .B1(_151_),
  .B2(_040_),
  .ZN(_041_)
);

NAND2_X1 _287_ (
  .A1(_029_),
  .A2(_130_),
  .ZN(_042_)
);

NOR2_X1 _288_ (
  .A1(_129_),
  .A2(x[0]),
  .ZN(_043_)
);

OAI21_X1 _289_ (
  .A(_041_),
  .B1(_042_),
  .B2(_043_),
  .ZN(_044_)
);

AOI21_X1 _290_ (
  .A(_032_),
  .B1(_039_),
  .B2(_044_),
  .ZN(_003_)
);

NAND3_X1 _291_ (
  .A1(_141_),
  .A2(_112_),
  .A3(_114_),
  .ZN(_045_)
);

NAND2_X1 _292_ (
  .A1(_036_),
  .A2(_045_),
  .ZN(_046_)
);

NAND3_X1 _293_ (
  .A1(_141_),
  .A2(_112_),
  .A3(_130_),
  .ZN(_047_)
);

NAND2_X1 _294_ (
  .A1(_041_),
  .A2(_047_),
  .ZN(_048_)
);

NAND3_X1 _295_ (
  .A1(_046_),
  .A2(_048_),
  .A3(_102_),
  .ZN(_049_)
);

NAND2_X1 _296_ (
  .A1(_103_),
  .A2(\coef[26] ),
  .ZN(_050_)
);

NAND2_X1 _297_ (
  .A1(_049_),
  .A2(_050_),
  .ZN(_004_)
);

NOR2_X1 _298_ (
  .A1(_102_),
  .A2(\coef[13] ),
  .ZN(_051_)
);

NAND3_X1 _299_ (
  .A1(_024_),
  .A2(_121_),
  .A3(_025_),
  .ZN(_052_)
);

INV_X1 _300_ (
  .A(_052_),
  .ZN(_053_)
);

OAI21_X1 _301_ (
  .A(_114_),
  .B1(_053_),
  .B2(_028_),
  .ZN(_054_)
);

INV_X1 _302_ (
  .A(_187_),
  .ZN(_055_)
);

NAND2_X1 _303_ (
  .A1(_106_),
  .A2(_055_),
  .ZN(_056_)
);

NAND2_X2 _304_ (
  .A1(_126_),
  .A2(_173_),
  .ZN(_057_)
);

NAND3_X1 _305_ (
  .A1(_056_),
  .A2(_109_),
  .A3(_057_),
  .ZN(_058_)
);

INV_X1 _306_ (
  .A(_058_),
  .ZN(_059_)
);

NOR2_X1 _307_ (
  .A1(_171_),
  .A2(_129_),
  .ZN(_060_)
);

OAI21_X1 _308_ (
  .A(_130_),
  .B1(_059_),
  .B2(_060_),
  .ZN(_061_)
);

NAND2_X1 _309_ (
  .A1(_054_),
  .A2(_061_),
  .ZN(_062_)
);

NAND2_X1 _310_ (
  .A1(_062_),
  .A2(_134_),
  .ZN(_063_)
);

NAND3_X1 _311_ (
  .A1(_017_),
  .A2(_018_),
  .A3(_129_),
  .ZN(_064_)
);

NAND2_X2 _312_ (
  .A1(_121_),
  .A2(_126_),
  .ZN(_065_)
);

NAND2_X1 _313_ (
  .A1(_065_),
  .A2(_113_),
  .ZN(_066_)
);

INV_X1 _314_ (
  .A(_066_),
  .ZN(_067_)
);

AOI21_X1 _315_ (
  .A(_134_),
  .B1(_064_),
  .B2(_067_),
  .ZN(_068_)
);

INV_X1 _316_ (
  .A(_185_),
  .ZN(_069_)
);

NAND2_X1 _317_ (
  .A1(_106_),
  .A2(_069_),
  .ZN(_070_)
);

NAND2_X1 _318_ (
  .A1(_126_),
  .A2(_175_),
  .ZN(_071_)
);

NAND3_X1 _319_ (
  .A1(_070_),
  .A2(_121_),
  .A3(_071_),
  .ZN(_072_)
);

NAND2_X1 _320_ (
  .A1(_072_),
  .A2(_037_),
  .ZN(_073_)
);

NAND2_X1 _321_ (
  .A1(_073_),
  .A2(_114_),
  .ZN(_074_)
);

AOI21_X1 _322_ (
  .A(_103_),
  .B1(_068_),
  .B2(_074_),
  .ZN(_075_)
);

AOI21_X2 _323_ (
  .A(_051_),
  .B1(_063_),
  .B2(_075_),
  .ZN(_005_)
);

NAND3_X1 _324_ (
  .A1(_070_),
  .A2(_109_),
  .A3(_071_),
  .ZN(_076_)
);

NAND2_X1 _325_ (
  .A1(_112_),
  .A2(_076_),
  .ZN(_077_)
);

NAND2_X1 _326_ (
  .A1(_077_),
  .A2(_130_),
  .ZN(_078_)
);

NAND3_X1 _327_ (
  .A1(_078_),
  .A2(_027_),
  .A3(_132_),
  .ZN(_079_)
);

NAND3_X1 _328_ (
  .A1(_138_),
  .A2(_129_),
  .A3(_139_),
  .ZN(_080_)
);

NAND3_X1 _329_ (
  .A1(_056_),
  .A2(_121_),
  .A3(_057_),
  .ZN(_081_)
);

NAND3_X1 _330_ (
  .A1(_080_),
  .A2(_081_),
  .A3(_114_),
  .ZN(_082_)
);

NAND3_X1 _331_ (
  .A1(_020_),
  .A2(_082_),
  .A3(_134_),
  .ZN(_083_)
);

NAND2_X1 _332_ (
  .A1(_079_),
  .A2(_083_),
  .ZN(_084_)
);

NAND2_X1 _333_ (
  .A1(_084_),
  .A2(_102_),
  .ZN(_085_)
);

NAND2_X1 _334_ (
  .A1(_103_),
  .A2(\coef[28] ),
  .ZN(_086_)
);

NAND2_X1 _335_ (
  .A1(_085_),
  .A2(_086_),
  .ZN(_006_)
);

NAND2_X1 _336_ (
  .A1(_010_),
  .A2(_029_),
  .ZN(_087_)
);

NAND2_X1 _337_ (
  .A1(_087_),
  .A2(_114_),
  .ZN(_088_)
);

NAND3_X1 _338_ (
  .A1(_118_),
  .A2(_119_),
  .A3(_129_),
  .ZN(_089_)
);

NAND3_X1 _339_ (
  .A1(_089_),
  .A2(_072_),
  .A3(_130_),
  .ZN(_090_)
);

NAND3_X1 _340_ (
  .A1(_088_),
  .A2(_090_),
  .A3(_132_),
  .ZN(_091_)
);

NAND3_X1 _341_ (
  .A1(_118_),
  .A2(_119_),
  .A3(_121_),
  .ZN(_092_)
);

NAND3_X1 _342_ (
  .A1(_092_),
  .A2(_058_),
  .A3(_114_),
  .ZN(_093_)
);

NAND3_X1 _343_ (
  .A1(_158_),
  .A2(_130_),
  .A3(_065_),
  .ZN(_094_)
);

NAND2_X1 _344_ (
  .A1(_093_),
  .A2(_094_),
  .ZN(_095_)
);

NAND2_X1 _345_ (
  .A1(_095_),
  .A2(_134_),
  .ZN(_096_)
);

NAND3_X1 _346_ (
  .A1(_091_),
  .A2(_096_),
  .A3(_102_),
  .ZN(_097_)
);

NAND2_X1 _347_ (
  .A1(_103_),
  .A2(\coef[29] ),
  .ZN(_098_)
);

NAND2_X1 _348_ (
  .A1(_097_),
  .A2(_098_),
  .ZN(_007_)
);

AOI21_X1 _349_ (
  .A(_103_),
  .B1(_149_),
  .B2(_134_),
  .ZN(_099_)
);

OAI21_X1 _350_ (
  .A(_099_),
  .B1(_134_),
  .B2(_128_),
  .ZN(_100_)
);

INV_X1 _351_ (
  .A(\coef[30] ),
  .ZN(_101_)
);

OAI21_X1 _352_ (
  .A(_100_),
  .B1(_102_),
  .B2(_101_),
  .ZN(_008_)
);

HA_X1 _353_ (
  .A(_171_),
  .B(_172_),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _354_ (
  .A(_171_),
  .B(_172_),
  .CO(_175_),
  .S(_176_)
);

HA_X1 _355_ (
  .A(_171_),
  .B(x[1]),
  .CO(_177_),
  .S(_178_)
);

HA_X1 _356_ (
  .A(_171_),
  .B(x[1]),
  .CO(_179_),
  .S(_180_)
);

HA_X1 _357_ (
  .A(x[0]),
  .B(_172_),
  .CO(_181_),
  .S(_182_)
);

HA_X1 _358_ (
  .A(x[0]),
  .B(_172_),
  .CO(_183_),
  .S(_184_)
);

HA_X1 _359_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_185_),
  .S(_186_)
);

HA_X1 _360_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_187_),
  .S(_188_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_170_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_169_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_168_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_167_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_166_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_165_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_164_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_163_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_162_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[28] , \coef[13] , \coef[26] , \coef[10] , \coef[24] , \coef[23] , \coef[10] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$e2471d3acfddfd8f107137e4952b02d9e7720f44\dctu

module \$paramod$e6bd937dcb54fb0697fee40c5f9824ba6fd53538\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire \coef[10] ;
wire \coef[11] ;
wire \coef[13] ;
wire \coef[15] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

BUF_X4 _30_ (
  .A(y[2]),
  .Z(_04_)
);

INV_X4 _31_ (
  .A(_04_),
  .ZN(_05_)
);

NAND2_X2 _32_ (
  .A1(_05_),
  .A2(y[1]),
  .ZN(_06_)
);

INV_X1 _33_ (
  .A(y[1]),
  .ZN(_07_)
);

NAND2_X1 _34_ (
  .A1(_07_),
  .A2(_04_),
  .ZN(_08_)
);

BUF_X4 _35_ (
  .A(ena),
  .Z(_09_)
);

NAND3_X1 _36_ (
  .A1(_06_),
  .A2(_08_),
  .A3(_09_),
  .ZN(_10_)
);

INV_X2 _37_ (
  .A(_09_),
  .ZN(_11_)
);

NAND2_X1 _38_ (
  .A1(_11_),
  .A2(\coef[11] ),
  .ZN(_12_)
);

NAND2_X1 _39_ (
  .A1(_10_),
  .A2(_12_),
  .ZN(_00_)
);

INV_X1 _40_ (
  .A(y[0]),
  .ZN(_13_)
);

NAND2_X2 _41_ (
  .A1(_05_),
  .A2(_13_),
  .ZN(_14_)
);

NAND2_X1 _42_ (
  .A1(_04_),
  .A2(y[0]),
  .ZN(_15_)
);

NAND3_X1 _43_ (
  .A1(_14_),
  .A2(_09_),
  .A3(_15_),
  .ZN(_16_)
);

NAND2_X1 _44_ (
  .A1(_11_),
  .A2(\coef[13] ),
  .ZN(_17_)
);

NAND2_X1 _45_ (
  .A1(_16_),
  .A2(_17_),
  .ZN(_01_)
);

NAND2_X1 _46_ (
  .A1(_13_),
  .A2(_04_),
  .ZN(_18_)
);

NAND2_X2 _47_ (
  .A1(_05_),
  .A2(y[0]),
  .ZN(_19_)
);

NAND3_X2 _48_ (
  .A1(_18_),
  .A2(_19_),
  .A3(_09_),
  .ZN(_20_)
);

NAND2_X1 _49_ (
  .A1(_11_),
  .A2(\coef[10] ),
  .ZN(_21_)
);

NAND2_X2 _50_ (
  .A1(_20_),
  .A2(_21_),
  .ZN(_02_)
);

NAND2_X1 _51_ (
  .A1(_11_),
  .A2(\coef[15] ),
  .ZN(_22_)
);

NAND2_X1 _52_ (
  .A1(_04_),
  .A2(y[1]),
  .ZN(_23_)
);

NAND2_X1 _53_ (
  .A1(_23_),
  .A2(_09_),
  .ZN(_24_)
);

NOR2_X1 _54_ (
  .A1(_04_),
  .A2(y[1]),
  .ZN(_25_)
);

OAI21_X2 _55_ (
  .A(_22_),
  .B1(_24_),
  .B2(_25_),
  .ZN(_03_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[11] ),
  .QN(_29_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_01_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_28_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_02_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_27_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_03_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_26_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[15] , \coef[15] , \coef[10] , \coef[13] , \coef[10] , \coef[15] , \coef[15] , \coef[11] , \coef[10] , \coef[11] , \coef[15] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$e6bd937dcb54fb0697fee40c5f9824ba6fd53538\dctu

module \$paramod$e9d96eb14c78f030ece167996f154f4849a68288\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _189_ (
  .A(x[1]),
  .ZN(_172_)
);

INV_X1 _190_ (
  .A(x[0]),
  .ZN(_171_)
);

BUF_X1 _191_ (
  .A(ena),
  .Z(_103_)
);

NOR2_X1 _192_ (
  .A1(\coef[21] ),
  .A2(_103_),
  .ZN(_104_)
);

INV_X2 _193_ (
  .A(x[2]),
  .ZN(_105_)
);

BUF_X8 _194_ (
  .A(_105_),
  .Z(_106_)
);

NAND2_X1 _195_ (
  .A1(_106_),
  .A2(_177_),
  .ZN(_107_)
);

INV_X1 _196_ (
  .A(_183_),
  .ZN(_108_)
);

BUF_X4 _197_ (
  .A(x[2]),
  .Z(_109_)
);

NAND2_X1 _198_ (
  .A1(_108_),
  .A2(_109_),
  .ZN(_110_)
);

BUF_X4 _199_ (
  .A(y[0]),
  .Z(_111_)
);

INV_X4 _200_ (
  .A(_111_),
  .ZN(_112_)
);

NAND3_X2 _201_ (
  .A1(_107_),
  .A2(_110_),
  .A3(_112_),
  .ZN(_113_)
);

INV_X1 _202_ (
  .A(_175_),
  .ZN(_114_)
);

NAND2_X2 _203_ (
  .A1(_106_),
  .A2(_114_),
  .ZN(_115_)
);

NAND2_X2 _204_ (
  .A1(_109_),
  .A2(_185_),
  .ZN(_116_)
);

NAND3_X1 _205_ (
  .A1(_115_),
  .A2(_111_),
  .A3(_116_),
  .ZN(_117_)
);

NAND2_X1 _206_ (
  .A1(_113_),
  .A2(_117_),
  .ZN(_118_)
);

BUF_X4 _207_ (
  .A(y[1]),
  .Z(_119_)
);

INV_X2 _208_ (
  .A(_119_),
  .ZN(_120_)
);

BUF_X4 _209_ (
  .A(y[2]),
  .Z(_121_)
);

NOR2_X2 _210_ (
  .A1(_120_),
  .A2(_121_),
  .ZN(_122_)
);

NAND2_X1 _211_ (
  .A1(_118_),
  .A2(_122_),
  .ZN(_123_)
);

NAND2_X2 _212_ (
  .A1(_106_),
  .A2(_179_),
  .ZN(_124_)
);

INV_X1 _213_ (
  .A(_181_),
  .ZN(_125_)
);

NAND2_X2 _214_ (
  .A1(_125_),
  .A2(_109_),
  .ZN(_126_)
);

BUF_X4 _215_ (
  .A(_111_),
  .Z(_127_)
);

NAND3_X1 _216_ (
  .A1(_124_),
  .A2(_126_),
  .A3(_127_),
  .ZN(_128_)
);

INV_X1 _217_ (
  .A(_173_),
  .ZN(_129_)
);

NAND2_X1 _218_ (
  .A1(_105_),
  .A2(_129_),
  .ZN(_130_)
);

NAND2_X4 _219_ (
  .A1(_109_),
  .A2(_187_),
  .ZN(_131_)
);

NAND3_X2 _220_ (
  .A1(_130_),
  .A2(_112_),
  .A3(_131_),
  .ZN(_132_)
);

NOR2_X1 _221_ (
  .A1(_119_),
  .A2(_121_),
  .ZN(_133_)
);

NAND3_X1 _222_ (
  .A1(_128_),
  .A2(_132_),
  .A3(_133_),
  .ZN(_134_)
);

NAND2_X1 _223_ (
  .A1(_123_),
  .A2(_134_),
  .ZN(_135_)
);

NAND2_X1 _224_ (
  .A1(_106_),
  .A2(_175_),
  .ZN(_136_)
);

INV_X1 _225_ (
  .A(_185_),
  .ZN(_137_)
);

NAND2_X1 _226_ (
  .A1(_137_),
  .A2(_109_),
  .ZN(_138_)
);

BUF_X8 _227_ (
  .A(_112_),
  .Z(_139_)
);

NAND3_X1 _228_ (
  .A1(_136_),
  .A2(_138_),
  .A3(_139_),
  .ZN(_140_)
);

INV_X1 _229_ (
  .A(_177_),
  .ZN(_141_)
);

NAND2_X1 _230_ (
  .A1(_106_),
  .A2(_141_),
  .ZN(_142_)
);

NAND2_X1 _231_ (
  .A1(_109_),
  .A2(_183_),
  .ZN(_143_)
);

NAND3_X1 _232_ (
  .A1(_142_),
  .A2(_111_),
  .A3(_143_),
  .ZN(_144_)
);

INV_X2 _233_ (
  .A(_121_),
  .ZN(_145_)
);

NOR2_X2 _234_ (
  .A1(_145_),
  .A2(_119_),
  .ZN(_146_)
);

AND3_X1 _235_ (
  .A1(_140_),
  .A2(_144_),
  .A3(_146_),
  .ZN(_147_)
);

NOR2_X2 _236_ (
  .A1(_135_),
  .A2(_147_),
  .ZN(_148_)
);

INV_X1 _237_ (
  .A(_103_),
  .ZN(_149_)
);

NAND3_X1 _238_ (
  .A1(_130_),
  .A2(_127_),
  .A3(_131_),
  .ZN(_150_)
);

NAND2_X1 _239_ (
  .A1(_119_),
  .A2(_121_),
  .ZN(_151_)
);

INV_X1 _240_ (
  .A(_151_),
  .ZN(_152_)
);

AND2_X1 _241_ (
  .A1(_150_),
  .A2(_152_),
  .ZN(_153_)
);

NAND3_X1 _242_ (
  .A1(_124_),
  .A2(_126_),
  .A3(_139_),
  .ZN(_154_)
);

AOI21_X1 _243_ (
  .A(_149_),
  .B1(_153_),
  .B2(_154_),
  .ZN(_155_)
);

AOI21_X2 _244_ (
  .A(_104_),
  .B1(_148_),
  .B2(_155_),
  .ZN(_000_)
);

NAND2_X1 _245_ (
  .A1(_105_),
  .A2(_183_),
  .ZN(_156_)
);

NAND2_X1 _246_ (
  .A1(_141_),
  .A2(x[2]),
  .ZN(_157_)
);

AND2_X1 _247_ (
  .A1(_156_),
  .A2(_157_),
  .ZN(_158_)
);

OAI21_X1 _248_ (
  .A(_158_),
  .B1(_122_),
  .B2(_146_),
  .ZN(_159_)
);

NOR2_X2 _249_ (
  .A1(_122_),
  .A2(_146_),
  .ZN(_160_)
);

NAND2_X2 _250_ (
  .A1(_109_),
  .A2(_179_),
  .ZN(_010_)
);

NAND2_X2 _251_ (
  .A1(_106_),
  .A2(_125_),
  .ZN(_011_)
);

NAND3_X1 _252_ (
  .A1(_160_),
  .A2(_010_),
  .A3(_011_),
  .ZN(_012_)
);

CLKBUF_X2 _253_ (
  .A(_103_),
  .Z(_013_)
);

NAND3_X1 _254_ (
  .A1(_159_),
  .A2(_012_),
  .A3(_013_),
  .ZN(_014_)
);

INV_X1 _255_ (
  .A(\coef[22] ),
  .ZN(_015_)
);

OAI21_X1 _256_ (
  .A(_014_),
  .B1(_013_),
  .B2(_015_),
  .ZN(_001_)
);

NOR2_X1 _257_ (
  .A1(_013_),
  .A2(\coef[23] ),
  .ZN(_016_)
);

OAI21_X1 _258_ (
  .A(_120_),
  .B1(_106_),
  .B2(_112_),
  .ZN(_017_)
);

INV_X1 _259_ (
  .A(_017_),
  .ZN(_018_)
);

NAND2_X1 _260_ (
  .A1(_154_),
  .A2(_018_),
  .ZN(_019_)
);

AOI21_X2 _261_ (
  .A(_120_),
  .B1(_139_),
  .B2(_106_),
  .ZN(_020_)
);

NAND2_X1 _262_ (
  .A1(_144_),
  .A2(_020_),
  .ZN(_021_)
);

NAND2_X1 _263_ (
  .A1(_019_),
  .A2(_021_),
  .ZN(_022_)
);

AOI21_X2 _264_ (
  .A(_149_),
  .B1(_022_),
  .B2(_145_),
  .ZN(_023_)
);

NAND2_X1 _265_ (
  .A1(_124_),
  .A2(_126_),
  .ZN(_024_)
);

NAND2_X1 _266_ (
  .A1(_024_),
  .A2(_127_),
  .ZN(_025_)
);

NAND2_X1 _267_ (
  .A1(_025_),
  .A2(_020_),
  .ZN(_026_)
);

NAND2_X1 _268_ (
  .A1(_113_),
  .A2(_018_),
  .ZN(_027_)
);

NAND3_X1 _269_ (
  .A1(_026_),
  .A2(_027_),
  .A3(_121_),
  .ZN(_028_)
);

AOI21_X2 _270_ (
  .A(_016_),
  .B1(_023_),
  .B2(_028_),
  .ZN(_002_)
);

NOR2_X1 _271_ (
  .A1(_013_),
  .A2(\coef[24] ),
  .ZN(_029_)
);

XNOR2_X1 _272_ (
  .A(_109_),
  .B(_174_),
  .ZN(_030_)
);

XNOR2_X1 _273_ (
  .A(_160_),
  .B(_030_),
  .ZN(_031_)
);

AOI21_X2 _274_ (
  .A(_029_),
  .B1(_031_),
  .B2(_013_),
  .ZN(_003_)
);

NOR2_X1 _275_ (
  .A1(_013_),
  .A2(\coef[25] ),
  .ZN(_032_)
);

NAND3_X2 _276_ (
  .A1(_115_),
  .A2(_139_),
  .A3(_116_),
  .ZN(_033_)
);

NAND2_X1 _277_ (
  .A1(x[1]),
  .A2(_127_),
  .ZN(_034_)
);

NAND2_X1 _278_ (
  .A1(_033_),
  .A2(_034_),
  .ZN(_035_)
);

NAND2_X1 _279_ (
  .A1(_035_),
  .A2(_146_),
  .ZN(_036_)
);

NAND2_X1 _280_ (
  .A1(_112_),
  .A2(x[1]),
  .ZN(_037_)
);

NAND3_X1 _281_ (
  .A1(_150_),
  .A2(_152_),
  .A3(_037_),
  .ZN(_038_)
);

NAND2_X1 _282_ (
  .A1(_036_),
  .A2(_038_),
  .ZN(_039_)
);

NAND3_X1 _283_ (
  .A1(_132_),
  .A2(_133_),
  .A3(_034_),
  .ZN(_040_)
);

INV_X1 _284_ (
  .A(_040_),
  .ZN(_041_)
);

NOR2_X2 _285_ (
  .A1(_039_),
  .A2(_041_),
  .ZN(_042_)
);

NAND2_X1 _286_ (
  .A1(_117_),
  .A2(_037_),
  .ZN(_043_)
);

AOI21_X1 _287_ (
  .A(_149_),
  .B1(_043_),
  .B2(_122_),
  .ZN(_044_)
);

AOI21_X2 _288_ (
  .A(_032_),
  .B1(_042_),
  .B2(_044_),
  .ZN(_004_)
);

NOR2_X1 _289_ (
  .A1(_013_),
  .A2(\coef[26] ),
  .ZN(_045_)
);

NAND2_X1 _290_ (
  .A1(_171_),
  .A2(_111_),
  .ZN(_046_)
);

NAND3_X1 _291_ (
  .A1(_046_),
  .A2(_119_),
  .A3(_145_),
  .ZN(_047_)
);

INV_X1 _292_ (
  .A(_047_),
  .ZN(_048_)
);

AOI21_X1 _293_ (
  .A(_149_),
  .B1(_048_),
  .B2(_132_),
  .ZN(_049_)
);

NAND3_X2 _294_ (
  .A1(_136_),
  .A2(_138_),
  .A3(_127_),
  .ZN(_050_)
);

AOI21_X2 _295_ (
  .A(_119_),
  .B1(_139_),
  .B2(x[0]),
  .ZN(_051_)
);

NAND3_X1 _296_ (
  .A1(_050_),
  .A2(_145_),
  .A3(_051_),
  .ZN(_052_)
);

AND2_X1 _297_ (
  .A1(_049_),
  .A2(_052_),
  .ZN(_053_)
);

NAND3_X1 _298_ (
  .A1(_033_),
  .A2(_119_),
  .A3(_046_),
  .ZN(_054_)
);

NAND2_X1 _299_ (
  .A1(_130_),
  .A2(_131_),
  .ZN(_055_)
);

NAND2_X1 _300_ (
  .A1(_055_),
  .A2(_127_),
  .ZN(_056_)
);

NAND2_X1 _301_ (
  .A1(_056_),
  .A2(_051_),
  .ZN(_057_)
);

NAND3_X1 _302_ (
  .A1(_054_),
  .A2(_121_),
  .A3(_057_),
  .ZN(_058_)
);

AOI21_X2 _303_ (
  .A(_045_),
  .B1(_053_),
  .B2(_058_),
  .ZN(_005_)
);

NOR2_X1 _304_ (
  .A1(_013_),
  .A2(\coef[27] ),
  .ZN(_059_)
);

NAND2_X1 _305_ (
  .A1(_106_),
  .A2(_187_),
  .ZN(_060_)
);

NAND2_X1 _306_ (
  .A1(_129_),
  .A2(_109_),
  .ZN(_061_)
);

NAND3_X1 _307_ (
  .A1(_060_),
  .A2(_061_),
  .A3(_139_),
  .ZN(_062_)
);

NAND3_X1 _308_ (
  .A1(_011_),
  .A2(_127_),
  .A3(_010_),
  .ZN(_063_)
);

NAND3_X1 _309_ (
  .A1(_062_),
  .A2(_063_),
  .A3(_122_),
  .ZN(_064_)
);

NAND2_X1 _310_ (
  .A1(_064_),
  .A2(_103_),
  .ZN(_065_)
);

NAND2_X1 _311_ (
  .A1(_158_),
  .A2(_139_),
  .ZN(_066_)
);

NAND2_X1 _312_ (
  .A1(_066_),
  .A2(_133_),
  .ZN(_067_)
);

NAND2_X1 _313_ (
  .A1(_106_),
  .A2(_137_),
  .ZN(_068_)
);

NAND2_X1 _314_ (
  .A1(_109_),
  .A2(_175_),
  .ZN(_069_)
);

NAND3_X1 _315_ (
  .A1(_068_),
  .A2(_127_),
  .A3(_069_),
  .ZN(_070_)
);

INV_X1 _316_ (
  .A(_070_),
  .ZN(_071_)
);

NOR2_X1 _317_ (
  .A1(_067_),
  .A2(_071_),
  .ZN(_072_)
);

NOR2_X1 _318_ (
  .A1(_065_),
  .A2(_072_),
  .ZN(_073_)
);

NAND3_X1 _319_ (
  .A1(_060_),
  .A2(_061_),
  .A3(_127_),
  .ZN(_074_)
);

NAND3_X1 _320_ (
  .A1(_011_),
  .A2(_139_),
  .A3(_010_),
  .ZN(_075_)
);

NAND3_X1 _321_ (
  .A1(_074_),
  .A2(_075_),
  .A3(_120_),
  .ZN(_076_)
);

NAND3_X1 _322_ (
  .A1(_156_),
  .A2(_157_),
  .A3(_127_),
  .ZN(_077_)
);

NAND3_X1 _323_ (
  .A1(_068_),
  .A2(_139_),
  .A3(_069_),
  .ZN(_078_)
);

NAND3_X1 _324_ (
  .A1(_077_),
  .A2(_078_),
  .A3(_119_),
  .ZN(_079_)
);

NAND2_X1 _325_ (
  .A1(_076_),
  .A2(_079_),
  .ZN(_080_)
);

NAND2_X1 _326_ (
  .A1(_080_),
  .A2(_121_),
  .ZN(_081_)
);

AOI21_X2 _327_ (
  .A(_059_),
  .B1(_073_),
  .B2(_081_),
  .ZN(_006_)
);

NOR2_X1 _328_ (
  .A1(_013_),
  .A2(\coef[28] ),
  .ZN(_082_)
);

NAND2_X1 _329_ (
  .A1(_025_),
  .A2(_113_),
  .ZN(_083_)
);

AOI21_X1 _330_ (
  .A(_149_),
  .B1(_083_),
  .B2(_145_),
  .ZN(_084_)
);

NAND3_X1 _331_ (
  .A1(_154_),
  .A2(_144_),
  .A3(_121_),
  .ZN(_085_)
);

AOI21_X1 _332_ (
  .A(_082_),
  .B1(_084_),
  .B2(_085_),
  .ZN(_007_)
);

NOR2_X1 _333_ (
  .A1(_013_),
  .A2(\coef[15] ),
  .ZN(_086_)
);

NAND2_X1 _334_ (
  .A1(_037_),
  .A2(_119_),
  .ZN(_087_)
);

INV_X1 _335_ (
  .A(_087_),
  .ZN(_088_)
);

NAND3_X1 _336_ (
  .A1(_050_),
  .A2(_145_),
  .A3(_088_),
  .ZN(_089_)
);

NAND2_X1 _337_ (
  .A1(_089_),
  .A2(_103_),
  .ZN(_090_)
);

NOR2_X1 _338_ (
  .A1(_139_),
  .A2(x[1]),
  .ZN(_091_)
);

INV_X1 _339_ (
  .A(_091_),
  .ZN(_092_)
);

NAND3_X1 _340_ (
  .A1(_132_),
  .A2(_133_),
  .A3(_092_),
  .ZN(_093_)
);

INV_X1 _341_ (
  .A(_093_),
  .ZN(_094_)
);

NOR2_X2 _342_ (
  .A1(_090_),
  .A2(_094_),
  .ZN(_095_)
);

AOI21_X1 _343_ (
  .A(_145_),
  .B1(_056_),
  .B2(_088_),
  .ZN(_096_)
);

NAND3_X1 _344_ (
  .A1(_033_),
  .A2(_120_),
  .A3(_092_),
  .ZN(_097_)
);

NAND2_X1 _345_ (
  .A1(_096_),
  .A2(_097_),
  .ZN(_098_)
);

AOI21_X2 _346_ (
  .A(_086_),
  .B1(_095_),
  .B2(_098_),
  .ZN(_008_)
);

NOR2_X1 _347_ (
  .A1(_103_),
  .A2(\coef[30] ),
  .ZN(_099_)
);

NAND3_X1 _348_ (
  .A1(_050_),
  .A2(_132_),
  .A3(_145_),
  .ZN(_100_)
);

AND2_X1 _349_ (
  .A1(_100_),
  .A2(_103_),
  .ZN(_101_)
);

NAND3_X1 _350_ (
  .A1(_140_),
  .A2(_150_),
  .A3(_121_),
  .ZN(_102_)
);

AOI21_X2 _351_ (
  .A(_099_),
  .B1(_101_),
  .B2(_102_),
  .ZN(_009_)
);

HA_X1 _352_ (
  .A(_171_),
  .B(_172_),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _353_ (
  .A(_171_),
  .B(_172_),
  .CO(_175_),
  .S(_176_)
);

HA_X1 _354_ (
  .A(_171_),
  .B(x[1]),
  .CO(_177_),
  .S(_178_)
);

HA_X1 _355_ (
  .A(_171_),
  .B(x[1]),
  .CO(_179_),
  .S(_180_)
);

HA_X1 _356_ (
  .A(x[0]),
  .B(_172_),
  .CO(_181_),
  .S(_182_)
);

HA_X1 _357_ (
  .A(x[0]),
  .B(_172_),
  .CO(_183_),
  .S(_184_)
);

HA_X1 _358_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_185_),
  .S(_186_)
);

HA_X1 _359_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_187_),
  .S(_188_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_170_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_169_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_168_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_167_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_166_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_165_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_164_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_163_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_162_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_161_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$e9d96eb14c78f030ece167996f154f4849a68288\dctu

module \$paramod$eb0441514cb1002bdcaf5201d3067d7bd1bbd3e9\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire \coef[10] ;
wire \coef[13] ;
wire \coef[29] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X2 _52_ (
  .A(x[2]),
  .ZN(_04_)
);

INV_X1 _53_ (
  .A(x[0]),
  .ZN(_05_)
);

NAND2_X1 _54_ (
  .A1(_04_),
  .A2(_05_),
  .ZN(_06_)
);

NAND2_X1 _55_ (
  .A1(x[2]),
  .A2(x[0]),
  .ZN(_07_)
);

NAND2_X1 _56_ (
  .A1(_06_),
  .A2(_07_),
  .ZN(_08_)
);

NAND2_X2 _57_ (
  .A1(_08_),
  .A2(y[0]),
  .ZN(_09_)
);

INV_X1 _58_ (
  .A(x[1]),
  .ZN(_10_)
);

NAND2_X1 _59_ (
  .A1(_04_),
  .A2(_10_),
  .ZN(_11_)
);

INV_X1 _60_ (
  .A(y[0]),
  .ZN(_12_)
);

NAND2_X1 _61_ (
  .A1(x[2]),
  .A2(x[1]),
  .ZN(_13_)
);

NAND3_X1 _62_ (
  .A1(_11_),
  .A2(_12_),
  .A3(_13_),
  .ZN(_14_)
);

NAND2_X1 _63_ (
  .A1(_09_),
  .A2(_14_),
  .ZN(_15_)
);

NAND2_X1 _64_ (
  .A1(_15_),
  .A2(y[1]),
  .ZN(_16_)
);

NAND2_X1 _65_ (
  .A1(_10_),
  .A2(x[2]),
  .ZN(_17_)
);

NAND2_X1 _66_ (
  .A1(_04_),
  .A2(x[1]),
  .ZN(_18_)
);

NAND3_X1 _67_ (
  .A1(_17_),
  .A2(_18_),
  .A3(y[0]),
  .ZN(_19_)
);

NAND3_X1 _68_ (
  .A1(_06_),
  .A2(_12_),
  .A3(_07_),
  .ZN(_20_)
);

NAND2_X1 _69_ (
  .A1(_19_),
  .A2(_20_),
  .ZN(_21_)
);

INV_X1 _70_ (
  .A(y[1]),
  .ZN(_22_)
);

NAND2_X1 _71_ (
  .A1(_21_),
  .A2(_22_),
  .ZN(_23_)
);

INV_X1 _72_ (
  .A(y[2]),
  .ZN(_24_)
);

NAND3_X1 _73_ (
  .A1(_16_),
  .A2(_23_),
  .A3(_24_),
  .ZN(_25_)
);

NAND3_X1 _74_ (
  .A1(_19_),
  .A2(_20_),
  .A3(_22_),
  .ZN(_26_)
);

NAND3_X1 _75_ (
  .A1(_09_),
  .A2(_14_),
  .A3(y[1]),
  .ZN(_27_)
);

NAND3_X1 _76_ (
  .A1(_26_),
  .A2(_27_),
  .A3(y[2]),
  .ZN(_28_)
);

NAND3_X1 _77_ (
  .A1(_25_),
  .A2(_28_),
  .A3(ena),
  .ZN(_29_)
);

INV_X1 _78_ (
  .A(ena),
  .ZN(_30_)
);

NAND2_X1 _79_ (
  .A1(_30_),
  .A2(\coef[13] ),
  .ZN(_31_)
);

NAND2_X1 _80_ (
  .A1(_29_),
  .A2(_31_),
  .ZN(_00_)
);

NAND3_X1 _81_ (
  .A1(_16_),
  .A2(_23_),
  .A3(y[2]),
  .ZN(_32_)
);

NAND3_X1 _82_ (
  .A1(_26_),
  .A2(_27_),
  .A3(_24_),
  .ZN(_33_)
);

NAND3_X1 _83_ (
  .A1(_32_),
  .A2(_33_),
  .A3(ena),
  .ZN(_34_)
);

NAND2_X1 _84_ (
  .A1(_30_),
  .A2(\coef[10] ),
  .ZN(_35_)
);

NAND2_X1 _85_ (
  .A1(_34_),
  .A2(_35_),
  .ZN(_01_)
);

NAND3_X1 _86_ (
  .A1(_17_),
  .A2(_18_),
  .A3(_12_),
  .ZN(_36_)
);

NAND3_X1 _87_ (
  .A1(_09_),
  .A2(_36_),
  .A3(_22_),
  .ZN(_37_)
);

NAND3_X1 _88_ (
  .A1(_11_),
  .A2(y[0]),
  .A3(_13_),
  .ZN(_38_)
);

NAND3_X1 _89_ (
  .A1(_38_),
  .A2(_20_),
  .A3(y[1]),
  .ZN(_39_)
);

NAND2_X1 _90_ (
  .A1(_37_),
  .A2(_39_),
  .ZN(_40_)
);

NAND2_X1 _91_ (
  .A1(_40_),
  .A2(y[2]),
  .ZN(_41_)
);

NAND3_X1 _92_ (
  .A1(_37_),
  .A2(_39_),
  .A3(_24_),
  .ZN(_42_)
);

NAND3_X1 _93_ (
  .A1(_41_),
  .A2(_42_),
  .A3(ena),
  .ZN(_43_)
);

NAND2_X1 _94_ (
  .A1(_30_),
  .A2(\coef[29] ),
  .ZN(_44_)
);

NAND2_X1 _95_ (
  .A1(_43_),
  .A2(_44_),
  .ZN(_02_)
);

NAND2_X1 _96_ (
  .A1(_30_),
  .A2(\coef[30] ),
  .ZN(_45_)
);

NAND2_X1 _97_ (
  .A1(_36_),
  .A2(_38_),
  .ZN(_46_)
);

XNOR2_X1 _98_ (
  .A(_46_),
  .B(_24_),
  .ZN(_47_)
);

OAI21_X1 _99_ (
  .A(_45_),
  .B1(_47_),
  .B2(_30_),
  .ZN(_03_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_51_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_01_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_50_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_02_),
  .CK(clk),
  .Q(\coef[29] ),
  .QN(_49_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_03_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_48_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[29] , \coef[10] , \coef[13] , \coef[10] , \coef[10] , \coef[13] , \coef[10] , \coef[13] , \coef[10] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$eb0441514cb1002bdcaf5201d3067d7bd1bbd3e9\dctu

module \$paramod$11fa2caec0040cf5bdd9aac167c50c8009d1fe68\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _189_ (
  .A(x[0]),
  .ZN(_171_)
);

INV_X1 _190_ (
  .A(x[1]),
  .ZN(_172_)
);

BUF_X1 _191_ (
  .A(ena),
  .Z(_103_)
);

NOR2_X1 _192_ (
  .A1(\coef[21] ),
  .A2(_103_),
  .ZN(_104_)
);

BUF_X4 _193_ (
  .A(x[2]),
  .Z(_105_)
);

INV_X4 _194_ (
  .A(_105_),
  .ZN(_106_)
);

BUF_X16 _195_ (
  .A(_106_),
  .Z(_107_)
);

NAND2_X2 _196_ (
  .A1(_107_),
  .A2(_181_),
  .ZN(_108_)
);

INV_X1 _197_ (
  .A(_179_),
  .ZN(_109_)
);

BUF_X8 _198_ (
  .A(_105_),
  .Z(_110_)
);

NAND2_X1 _199_ (
  .A1(_109_),
  .A2(_110_),
  .ZN(_111_)
);

BUF_X4 _200_ (
  .A(y[0]),
  .Z(_112_)
);

NAND3_X2 _201_ (
  .A1(_108_),
  .A2(_111_),
  .A3(_112_),
  .ZN(_113_)
);

INV_X1 _202_ (
  .A(_187_),
  .ZN(_114_)
);

NAND2_X4 _203_ (
  .A1(_107_),
  .A2(_114_),
  .ZN(_115_)
);

INV_X4 _204_ (
  .A(_112_),
  .ZN(_116_)
);

NAND2_X1 _205_ (
  .A1(_105_),
  .A2(_173_),
  .ZN(_117_)
);

NAND3_X4 _206_ (
  .A1(_115_),
  .A2(_116_),
  .A3(_117_),
  .ZN(_118_)
);

NAND2_X1 _207_ (
  .A1(_113_),
  .A2(_118_),
  .ZN(_119_)
);

BUF_X4 _208_ (
  .A(y[2]),
  .Z(_120_)
);

INV_X4 _209_ (
  .A(_120_),
  .ZN(_121_)
);

BUF_X4 _210_ (
  .A(y[1]),
  .Z(_122_)
);

NAND2_X1 _211_ (
  .A1(_121_),
  .A2(_122_),
  .ZN(_123_)
);

INV_X1 _212_ (
  .A(_123_),
  .ZN(_124_)
);

NAND2_X1 _213_ (
  .A1(_119_),
  .A2(_124_),
  .ZN(_125_)
);

NAND2_X4 _214_ (
  .A1(_115_),
  .A2(_117_),
  .ZN(_126_)
);

BUF_X4 _215_ (
  .A(_112_),
  .Z(_127_)
);

NAND2_X2 _216_ (
  .A1(_126_),
  .A2(_127_),
  .ZN(_128_)
);

INV_X1 _217_ (
  .A(_181_),
  .ZN(_129_)
);

NAND2_X4 _218_ (
  .A1(_107_),
  .A2(_129_),
  .ZN(_130_)
);

BUF_X8 _219_ (
  .A(_116_),
  .Z(_131_)
);

NAND2_X2 _220_ (
  .A1(_110_),
  .A2(_179_),
  .ZN(_132_)
);

NAND3_X2 _221_ (
  .A1(_130_),
  .A2(_131_),
  .A3(_132_),
  .ZN(_133_)
);

NOR2_X4 _222_ (
  .A1(_121_),
  .A2(_122_),
  .ZN(_134_)
);

NAND3_X1 _223_ (
  .A1(_128_),
  .A2(_133_),
  .A3(_134_),
  .ZN(_135_)
);

NAND2_X1 _224_ (
  .A1(_125_),
  .A2(_135_),
  .ZN(_136_)
);

NOR2_X1 _225_ (
  .A1(_122_),
  .A2(_120_),
  .ZN(_137_)
);

INV_X1 _226_ (
  .A(_137_),
  .ZN(_138_)
);

INV_X1 _227_ (
  .A(_185_),
  .ZN(_139_)
);

NAND2_X4 _228_ (
  .A1(_107_),
  .A2(_139_),
  .ZN(_140_)
);

NAND2_X1 _229_ (
  .A1(_110_),
  .A2(_175_),
  .ZN(_141_)
);

NAND2_X1 _230_ (
  .A1(_140_),
  .A2(_141_),
  .ZN(_142_)
);

NAND2_X2 _231_ (
  .A1(_142_),
  .A2(_127_),
  .ZN(_143_)
);

INV_X1 _232_ (
  .A(_183_),
  .ZN(_144_)
);

NAND2_X2 _233_ (
  .A1(_107_),
  .A2(_144_),
  .ZN(_145_)
);

NAND2_X1 _234_ (
  .A1(_105_),
  .A2(_177_),
  .ZN(_146_)
);

NAND3_X1 _235_ (
  .A1(_145_),
  .A2(_131_),
  .A3(_146_),
  .ZN(_147_)
);

AOI21_X1 _236_ (
  .A(_138_),
  .B1(_143_),
  .B2(_147_),
  .ZN(_148_)
);

NOR2_X2 _237_ (
  .A1(_136_),
  .A2(_148_),
  .ZN(_149_)
);

INV_X1 _238_ (
  .A(_103_),
  .ZN(_150_)
);

NAND2_X4 _239_ (
  .A1(_107_),
  .A2(_183_),
  .ZN(_151_)
);

INV_X1 _240_ (
  .A(_177_),
  .ZN(_152_)
);

NAND2_X2 _241_ (
  .A1(_152_),
  .A2(_110_),
  .ZN(_153_)
);

NAND3_X1 _242_ (
  .A1(_151_),
  .A2(_153_),
  .A3(_127_),
  .ZN(_154_)
);

NAND2_X1 _243_ (
  .A1(_122_),
  .A2(_120_),
  .ZN(_155_)
);

INV_X1 _244_ (
  .A(_155_),
  .ZN(_156_)
);

AND2_X1 _245_ (
  .A1(_154_),
  .A2(_156_),
  .ZN(_157_)
);

NAND3_X1 _246_ (
  .A1(_140_),
  .A2(_131_),
  .A3(_141_),
  .ZN(_158_)
);

AOI21_X1 _247_ (
  .A(_150_),
  .B1(_157_),
  .B2(_158_),
  .ZN(_159_)
);

AOI21_X2 _248_ (
  .A(_104_),
  .B1(_149_),
  .B2(_159_),
  .ZN(_000_)
);

INV_X1 _249_ (
  .A(_134_),
  .ZN(_160_)
);

NAND2_X1 _250_ (
  .A1(_160_),
  .A2(_123_),
  .ZN(_010_)
);

NAND2_X1 _251_ (
  .A1(_107_),
  .A2(_175_),
  .ZN(_011_)
);

NAND2_X1 _252_ (
  .A1(_139_),
  .A2(_110_),
  .ZN(_012_)
);

NAND3_X1 _253_ (
  .A1(_010_),
  .A2(_011_),
  .A3(_012_),
  .ZN(_013_)
);

INV_X1 _254_ (
  .A(_173_),
  .ZN(_014_)
);

NAND2_X1 _255_ (
  .A1(_107_),
  .A2(_014_),
  .ZN(_015_)
);

NAND2_X1 _256_ (
  .A1(_110_),
  .A2(_187_),
  .ZN(_016_)
);

NAND4_X1 _257_ (
  .A1(_160_),
  .A2(_015_),
  .A3(_123_),
  .A4(_016_),
  .ZN(_017_)
);

BUF_X1 _258_ (
  .A(_103_),
  .Z(_018_)
);

NAND3_X1 _259_ (
  .A1(_013_),
  .A2(_017_),
  .A3(_018_),
  .ZN(_019_)
);

INV_X1 _260_ (
  .A(\coef[22] ),
  .ZN(_020_)
);

OAI21_X1 _261_ (
  .A(_019_),
  .B1(_018_),
  .B2(_020_),
  .ZN(_001_)
);

NOR2_X1 _262_ (
  .A1(_018_),
  .A2(\coef[23] ),
  .ZN(_021_)
);

OAI21_X1 _263_ (
  .A(_122_),
  .B1(_171_),
  .B2(_112_),
  .ZN(_022_)
);

INV_X1 _264_ (
  .A(_022_),
  .ZN(_023_)
);

NAND2_X1 _265_ (
  .A1(_128_),
  .A2(_023_),
  .ZN(_024_)
);

AOI21_X1 _266_ (
  .A(_122_),
  .B1(_171_),
  .B2(_112_),
  .ZN(_025_)
);

NAND2_X1 _267_ (
  .A1(_158_),
  .A2(_025_),
  .ZN(_026_)
);

NAND2_X1 _268_ (
  .A1(_024_),
  .A2(_026_),
  .ZN(_027_)
);

AOI21_X2 _269_ (
  .A(_150_),
  .B1(_027_),
  .B2(_121_),
  .ZN(_028_)
);

NAND2_X1 _270_ (
  .A1(_143_),
  .A2(_023_),
  .ZN(_029_)
);

NAND2_X1 _271_ (
  .A1(_118_),
  .A2(_025_),
  .ZN(_030_)
);

NAND3_X1 _272_ (
  .A1(_029_),
  .A2(_030_),
  .A3(_120_),
  .ZN(_031_)
);

AOI21_X2 _273_ (
  .A(_021_),
  .B1(_028_),
  .B2(_031_),
  .ZN(_002_)
);

NOR2_X1 _274_ (
  .A1(_018_),
  .A2(\coef[24] ),
  .ZN(_032_)
);

XNOR2_X1 _275_ (
  .A(_010_),
  .B(_172_),
  .ZN(_033_)
);

AOI21_X1 _276_ (
  .A(_032_),
  .B1(_033_),
  .B2(_018_),
  .ZN(_003_)
);

NOR2_X1 _277_ (
  .A1(_018_),
  .A2(\coef[25] ),
  .ZN(_034_)
);

INV_X1 _278_ (
  .A(_174_),
  .ZN(_035_)
);

NAND2_X2 _279_ (
  .A1(_106_),
  .A2(_035_),
  .ZN(_036_)
);

NAND2_X1 _280_ (
  .A1(_105_),
  .A2(_174_),
  .ZN(_037_)
);

NAND2_X1 _281_ (
  .A1(_036_),
  .A2(_037_),
  .ZN(_038_)
);

NAND2_X1 _282_ (
  .A1(_038_),
  .A2(_127_),
  .ZN(_039_)
);

NAND3_X1 _283_ (
  .A1(_039_),
  .A2(_133_),
  .A3(_134_),
  .ZN(_040_)
);

NAND3_X1 _284_ (
  .A1(_036_),
  .A2(_116_),
  .A3(_037_),
  .ZN(_041_)
);

NAND3_X1 _285_ (
  .A1(_154_),
  .A2(_041_),
  .A3(_156_),
  .ZN(_042_)
);

NAND2_X1 _286_ (
  .A1(_040_),
  .A2(_042_),
  .ZN(_043_)
);

AOI21_X1 _287_ (
  .A(_138_),
  .B1(_039_),
  .B2(_147_),
  .ZN(_044_)
);

NOR2_X1 _288_ (
  .A1(_043_),
  .A2(_044_),
  .ZN(_045_)
);

NAND2_X1 _289_ (
  .A1(_113_),
  .A2(_041_),
  .ZN(_046_)
);

AOI21_X1 _290_ (
  .A(_150_),
  .B1(_046_),
  .B2(_124_),
  .ZN(_047_)
);

AOI21_X2 _291_ (
  .A(_034_),
  .B1(_045_),
  .B2(_047_),
  .ZN(_004_)
);

NOR2_X1 _292_ (
  .A1(_018_),
  .A2(\coef[26] ),
  .ZN(_048_)
);

NAND3_X2 _293_ (
  .A1(_151_),
  .A2(_153_),
  .A3(_131_),
  .ZN(_049_)
);

OAI21_X1 _294_ (
  .A(_122_),
  .B1(_116_),
  .B2(_110_),
  .ZN(_050_)
);

INV_X1 _295_ (
  .A(_050_),
  .ZN(_051_)
);

NAND2_X1 _296_ (
  .A1(_049_),
  .A2(_051_),
  .ZN(_052_)
);

NAND3_X2 _297_ (
  .A1(_130_),
  .A2(_127_),
  .A3(_132_),
  .ZN(_053_)
);

AOI21_X2 _298_ (
  .A(_122_),
  .B1(_131_),
  .B2(_110_),
  .ZN(_054_)
);

NAND2_X1 _299_ (
  .A1(_053_),
  .A2(_054_),
  .ZN(_055_)
);

NAND2_X1 _300_ (
  .A1(_052_),
  .A2(_055_),
  .ZN(_056_)
);

AOI21_X2 _301_ (
  .A(_150_),
  .B1(_056_),
  .B2(_121_),
  .ZN(_057_)
);

NAND3_X1 _302_ (
  .A1(_108_),
  .A2(_111_),
  .A3(_131_),
  .ZN(_058_)
);

NAND2_X1 _303_ (
  .A1(_058_),
  .A2(_051_),
  .ZN(_059_)
);

NAND3_X2 _304_ (
  .A1(_145_),
  .A2(_112_),
  .A3(_146_),
  .ZN(_060_)
);

NAND2_X1 _305_ (
  .A1(_060_),
  .A2(_054_),
  .ZN(_061_)
);

NAND3_X1 _306_ (
  .A1(_059_),
  .A2(_061_),
  .A3(_120_),
  .ZN(_062_)
);

AOI21_X2 _307_ (
  .A(_048_),
  .B1(_057_),
  .B2(_062_),
  .ZN(_005_)
);

NOR2_X1 _308_ (
  .A1(_018_),
  .A2(\coef[27] ),
  .ZN(_063_)
);

NAND3_X1 _309_ (
  .A1(_011_),
  .A2(_012_),
  .A3(_127_),
  .ZN(_064_)
);

NAND2_X1 _310_ (
  .A1(_107_),
  .A2(_152_),
  .ZN(_065_)
);

NAND2_X1 _311_ (
  .A1(_110_),
  .A2(_183_),
  .ZN(_066_)
);

NAND3_X1 _312_ (
  .A1(_065_),
  .A2(_131_),
  .A3(_066_),
  .ZN(_067_)
);

NAND3_X1 _313_ (
  .A1(_064_),
  .A2(_067_),
  .A3(_156_),
  .ZN(_068_)
);

NAND3_X1 _314_ (
  .A1(_011_),
  .A2(_012_),
  .A3(_131_),
  .ZN(_069_)
);

NAND3_X1 _315_ (
  .A1(_065_),
  .A2(_127_),
  .A3(_066_),
  .ZN(_070_)
);

NAND3_X1 _316_ (
  .A1(_069_),
  .A2(_070_),
  .A3(_137_),
  .ZN(_071_)
);

NAND2_X1 _317_ (
  .A1(_068_),
  .A2(_071_),
  .ZN(_072_)
);

NAND2_X1 _318_ (
  .A1(_107_),
  .A2(_109_),
  .ZN(_073_)
);

NAND2_X1 _319_ (
  .A1(_110_),
  .A2(_181_),
  .ZN(_074_)
);

NAND2_X1 _320_ (
  .A1(_073_),
  .A2(_074_),
  .ZN(_075_)
);

NAND2_X1 _321_ (
  .A1(_075_),
  .A2(_127_),
  .ZN(_076_)
);

NAND3_X1 _322_ (
  .A1(_015_),
  .A2(_131_),
  .A3(_016_),
  .ZN(_077_)
);

AND3_X2 _323_ (
  .A1(_076_),
  .A2(_077_),
  .A3(_134_),
  .ZN(_078_)
);

NOR2_X2 _324_ (
  .A1(_072_),
  .A2(_078_),
  .ZN(_079_)
);

NAND2_X1 _325_ (
  .A1(_075_),
  .A2(_131_),
  .ZN(_080_)
);

NAND3_X1 _326_ (
  .A1(_015_),
  .A2(_127_),
  .A3(_016_),
  .ZN(_081_)
);

NAND3_X1 _327_ (
  .A1(_080_),
  .A2(_081_),
  .A3(_124_),
  .ZN(_082_)
);

NAND2_X1 _328_ (
  .A1(_082_),
  .A2(_103_),
  .ZN(_083_)
);

INV_X1 _329_ (
  .A(_083_),
  .ZN(_084_)
);

AOI21_X2 _330_ (
  .A(_063_),
  .B1(_079_),
  .B2(_084_),
  .ZN(_006_)
);

NOR2_X1 _331_ (
  .A1(_018_),
  .A2(\coef[28] ),
  .ZN(_085_)
);

NAND2_X1 _332_ (
  .A1(_143_),
  .A2(_118_),
  .ZN(_086_)
);

AOI21_X1 _333_ (
  .A(_150_),
  .B1(_086_),
  .B2(_121_),
  .ZN(_087_)
);

NAND3_X1 _334_ (
  .A1(_128_),
  .A2(_158_),
  .A3(_120_),
  .ZN(_088_)
);

AOI21_X1 _335_ (
  .A(_085_),
  .B1(_087_),
  .B2(_088_),
  .ZN(_007_)
);

NAND2_X1 _336_ (
  .A1(_060_),
  .A2(_041_),
  .ZN(_089_)
);

NAND2_X1 _337_ (
  .A1(_089_),
  .A2(_156_),
  .ZN(_090_)
);

NAND3_X1 _338_ (
  .A1(_036_),
  .A2(_127_),
  .A3(_037_),
  .ZN(_091_)
);

NAND3_X1 _339_ (
  .A1(_133_),
  .A2(_091_),
  .A3(_134_),
  .ZN(_092_)
);

NAND3_X1 _340_ (
  .A1(_090_),
  .A2(_092_),
  .A3(_103_),
  .ZN(_093_)
);

NAND3_X1 _341_ (
  .A1(_039_),
  .A2(_049_),
  .A3(_137_),
  .ZN(_094_)
);

NAND3_X1 _342_ (
  .A1(_053_),
  .A2(_041_),
  .A3(_124_),
  .ZN(_095_)
);

NAND2_X1 _343_ (
  .A1(_094_),
  .A2(_095_),
  .ZN(_096_)
);

NOR2_X2 _344_ (
  .A1(_093_),
  .A2(_096_),
  .ZN(_097_)
);

NOR2_X1 _345_ (
  .A1(_018_),
  .A2(\coef[15] ),
  .ZN(_098_)
);

NOR2_X2 _346_ (
  .A1(_097_),
  .A2(_098_),
  .ZN(_008_)
);

NOR2_X1 _347_ (
  .A1(_103_),
  .A2(\coef[30] ),
  .ZN(_099_)
);

NAND2_X1 _348_ (
  .A1(_058_),
  .A2(_060_),
  .ZN(_100_)
);

AOI21_X1 _349_ (
  .A(_150_),
  .B1(_100_),
  .B2(_120_),
  .ZN(_101_)
);

NAND3_X1 _350_ (
  .A1(_049_),
  .A2(_053_),
  .A3(_121_),
  .ZN(_102_)
);

AOI21_X1 _351_ (
  .A(_099_),
  .B1(_101_),
  .B2(_102_),
  .ZN(_009_)
);

HA_X1 _352_ (
  .A(_171_),
  .B(_172_),
  .CO(_173_),
  .S(_174_)
);

HA_X1 _353_ (
  .A(_171_),
  .B(_172_),
  .CO(_175_),
  .S(_176_)
);

HA_X1 _354_ (
  .A(_171_),
  .B(x[1]),
  .CO(_177_),
  .S(_178_)
);

HA_X1 _355_ (
  .A(_171_),
  .B(x[1]),
  .CO(_179_),
  .S(_180_)
);

HA_X1 _356_ (
  .A(x[0]),
  .B(_172_),
  .CO(_181_),
  .S(_182_)
);

HA_X1 _357_ (
  .A(x[0]),
  .B(_172_),
  .CO(_183_),
  .S(_184_)
);

HA_X1 _358_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_185_),
  .S(_186_)
);

HA_X1 _359_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_187_),
  .S(_188_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_170_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_169_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_168_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_167_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_166_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_165_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_164_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_163_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_162_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_161_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$11fa2caec0040cf5bdd9aac167c50c8009d1fe68\dctu

module \$paramod$f06914ec453560c29e1738d8a2be788b84af024b\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire \coef[10] ;
wire \coef[11] ;
wire \coef[13] ;
wire \coef[15] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X2 _37_ (
  .A(x[2]),
  .ZN(_04_)
);

XNOR2_X1 _38_ (
  .A(_04_),
  .B(x[1]),
  .ZN(_05_)
);

INV_X1 _39_ (
  .A(y[0]),
  .ZN(_06_)
);

NAND2_X1 _40_ (
  .A1(_06_),
  .A2(y[1]),
  .ZN(_07_)
);

INV_X2 _41_ (
  .A(y[1]),
  .ZN(_08_)
);

NAND2_X1 _42_ (
  .A1(_08_),
  .A2(y[0]),
  .ZN(_09_)
);

NAND2_X1 _43_ (
  .A1(_07_),
  .A2(_09_),
  .ZN(_10_)
);

INV_X1 _44_ (
  .A(_10_),
  .ZN(_11_)
);

NAND2_X1 _45_ (
  .A1(_05_),
  .A2(_11_),
  .ZN(_12_)
);

XNOR2_X1 _46_ (
  .A(x[1]),
  .B(x[2]),
  .ZN(_13_)
);

NAND2_X1 _47_ (
  .A1(_13_),
  .A2(_10_),
  .ZN(_14_)
);

NAND3_X1 _48_ (
  .A1(_12_),
  .A2(_14_),
  .A3(ena),
  .ZN(_15_)
);

INV_X1 _49_ (
  .A(ena),
  .ZN(_16_)
);

NAND2_X1 _50_ (
  .A1(_16_),
  .A2(\coef[11] ),
  .ZN(_17_)
);

NAND2_X1 _51_ (
  .A1(_15_),
  .A2(_17_),
  .ZN(_00_)
);

NOR2_X1 _52_ (
  .A1(ena),
  .A2(\coef[13] ),
  .ZN(_18_)
);

NAND2_X2 _53_ (
  .A1(_08_),
  .A2(x[0]),
  .ZN(_19_)
);

INV_X1 _54_ (
  .A(x[0]),
  .ZN(_20_)
);

NAND2_X1 _55_ (
  .A1(_20_),
  .A2(y[1]),
  .ZN(_21_)
);

NAND2_X2 _56_ (
  .A1(_19_),
  .A2(_21_),
  .ZN(_22_)
);

NAND2_X1 _57_ (
  .A1(_04_),
  .A2(_06_),
  .ZN(_23_)
);

NAND2_X1 _58_ (
  .A1(x[2]),
  .A2(y[0]),
  .ZN(_24_)
);

NAND2_X2 _59_ (
  .A1(_23_),
  .A2(_24_),
  .ZN(_25_)
);

AOI21_X4 _60_ (
  .A(_16_),
  .B1(_22_),
  .B2(_25_),
  .ZN(_26_)
);

OR2_X4 _61_ (
  .A1(_25_),
  .A2(_22_),
  .ZN(_27_)
);

AOI21_X4 _62_ (
  .A(_18_),
  .B1(_26_),
  .B2(_27_),
  .ZN(_01_)
);

NAND2_X2 _63_ (
  .A1(_26_),
  .A2(_27_),
  .ZN(_28_)
);

NAND2_X1 _64_ (
  .A1(_16_),
  .A2(\coef[10] ),
  .ZN(_29_)
);

NAND2_X2 _65_ (
  .A1(_28_),
  .A2(_29_),
  .ZN(_02_)
);

NAND2_X1 _66_ (
  .A1(_12_),
  .A2(_14_),
  .ZN(_30_)
);

NAND2_X1 _67_ (
  .A1(_30_),
  .A2(ena),
  .ZN(_31_)
);

NAND2_X1 _68_ (
  .A1(_16_),
  .A2(\coef[15] ),
  .ZN(_32_)
);

NAND2_X1 _69_ (
  .A1(_31_),
  .A2(_32_),
  .ZN(_03_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[11] ),
  .QN(_36_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_01_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_35_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_02_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_34_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_03_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_33_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[15] , \coef[15] , \coef[10] , \coef[13] , \coef[10] , \coef[15] , \coef[15] , \coef[11] , \coef[10] , \coef[11] , \coef[15] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$f06914ec453560c29e1738d8a2be788b84af024b\dctu

module \$paramod$f1b01728a98736f8d413a71bd9a7600c5a6961e3\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _063_ (
  .A(y[0]),
  .ZN(_049_)
);

INV_X1 _064_ (
  .A(y[1]),
  .ZN(_050_)
);

INV_X1 _065_ (
  .A(_052_),
  .ZN(_008_)
);

BUF_X4 _066_ (
  .A(y[2]),
  .Z(_009_)
);

NAND2_X1 _067_ (
  .A1(_008_),
  .A2(_009_),
  .ZN(_010_)
);

INV_X4 _068_ (
  .A(_009_),
  .ZN(_011_)
);

NAND2_X2 _069_ (
  .A1(_011_),
  .A2(_052_),
  .ZN(_012_)
);

BUF_X4 _070_ (
  .A(ena),
  .Z(_013_)
);

NAND3_X1 _071_ (
  .A1(_010_),
  .A2(_012_),
  .A3(_013_),
  .ZN(_014_)
);

INV_X4 _072_ (
  .A(_013_),
  .ZN(_015_)
);

NAND2_X1 _073_ (
  .A1(_015_),
  .A2(\coef[21] ),
  .ZN(_016_)
);

NAND2_X1 _074_ (
  .A1(_014_),
  .A2(_016_),
  .ZN(_000_)
);

NAND2_X1 _075_ (
  .A1(_015_),
  .A2(\coef[22] ),
  .ZN(_017_)
);

NAND2_X1 _076_ (
  .A1(_009_),
  .A2(_057_),
  .ZN(_018_)
);

NAND2_X1 _077_ (
  .A1(_018_),
  .A2(_013_),
  .ZN(_019_)
);

NOR2_X1 _078_ (
  .A1(_009_),
  .A2(_055_),
  .ZN(_020_)
);

OAI21_X1 _079_ (
  .A(_017_),
  .B1(_019_),
  .B2(_020_),
  .ZN(_001_)
);

INV_X1 _080_ (
  .A(_061_),
  .ZN(_021_)
);

NAND2_X1 _081_ (
  .A1(_021_),
  .A2(_009_),
  .ZN(_022_)
);

NAND2_X2 _082_ (
  .A1(_011_),
  .A2(_051_),
  .ZN(_023_)
);

NAND3_X1 _083_ (
  .A1(_022_),
  .A2(_023_),
  .A3(_013_),
  .ZN(_024_)
);

NAND2_X1 _084_ (
  .A1(_015_),
  .A2(\coef[23] ),
  .ZN(_025_)
);

NAND2_X1 _085_ (
  .A1(_024_),
  .A2(_025_),
  .ZN(_002_)
);

INV_X1 _086_ (
  .A(_059_),
  .ZN(_026_)
);

NAND2_X1 _087_ (
  .A1(_026_),
  .A2(_009_),
  .ZN(_027_)
);

NAND2_X2 _088_ (
  .A1(_011_),
  .A2(_053_),
  .ZN(_028_)
);

NAND3_X1 _089_ (
  .A1(_027_),
  .A2(_028_),
  .A3(_013_),
  .ZN(_029_)
);

NAND2_X1 _090_ (
  .A1(_015_),
  .A2(\coef[14] ),
  .ZN(_030_)
);

NAND2_X1 _091_ (
  .A1(_029_),
  .A2(_030_),
  .ZN(_003_)
);

NAND2_X1 _092_ (
  .A1(_015_),
  .A2(\coef[13] ),
  .ZN(_031_)
);

OAI21_X1 _093_ (
  .A(_031_),
  .B1(y[0]),
  .B2(_015_),
  .ZN(_004_)
);

NAND2_X1 _094_ (
  .A1(_015_),
  .A2(\coef[28] ),
  .ZN(_032_)
);

OAI21_X1 _095_ (
  .A(_032_),
  .B1(y[1]),
  .B2(_015_),
  .ZN(_005_)
);

NAND2_X1 _096_ (
  .A1(_015_),
  .A2(\coef[15] ),
  .ZN(_033_)
);

NAND2_X1 _097_ (
  .A1(_009_),
  .A2(_051_),
  .ZN(_034_)
);

NAND2_X1 _098_ (
  .A1(_034_),
  .A2(_013_),
  .ZN(_035_)
);

NOR2_X1 _099_ (
  .A1(_009_),
  .A2(_061_),
  .ZN(_036_)
);

OAI21_X1 _100_ (
  .A(_033_),
  .B1(_035_),
  .B2(_036_),
  .ZN(_006_)
);

NAND2_X1 _101_ (
  .A1(_015_),
  .A2(\coef[12] ),
  .ZN(_037_)
);

NAND2_X1 _102_ (
  .A1(_009_),
  .A2(_053_),
  .ZN(_038_)
);

NAND2_X1 _103_ (
  .A1(_038_),
  .A2(_013_),
  .ZN(_039_)
);

NOR2_X1 _104_ (
  .A1(_009_),
  .A2(_059_),
  .ZN(_040_)
);

OAI21_X1 _105_ (
  .A(_037_),
  .B1(_039_),
  .B2(_040_),
  .ZN(_007_)
);

HA_X1 _106_ (
  .A(_049_),
  .B(_050_),
  .CO(_051_),
  .S(_052_)
);

HA_X1 _107_ (
  .A(_049_),
  .B(y[1]),
  .CO(_053_),
  .S(_054_)
);

HA_X1 _108_ (
  .A(_049_),
  .B(y[1]),
  .CO(_055_),
  .S(_056_)
);

HA_X1 _109_ (
  .A(y[0]),
  .B(_050_),
  .CO(_057_),
  .S(_058_)
);

HA_X1 _110_ (
  .A(y[0]),
  .B(_050_),
  .CO(_059_),
  .S(_060_)
);

HA_X1 _111_ (
  .A(y[0]),
  .B(y[1]),
  .CO(_061_),
  .S(_062_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_048_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_047_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_046_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_045_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_044_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_043_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_042_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_041_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$f1b01728a98736f8d413a71bd9a7600c5a6961e3\dctu

module \$paramod$f5bb6813249a03e2893277297591ec050ac518dc\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[24] ;
wire \coef[25] ;
wire \coef[26] ;
wire \coef[27] ;
wire \coef[28] ;
wire \coef[30] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

BUF_X2 _103_ (
  .A(y[2]),
  .Z(_027_)
);

INV_X2 _104_ (
  .A(_027_),
  .ZN(_028_)
);

INV_X2 _105_ (
  .A(x[2]),
  .ZN(_029_)
);

INV_X1 _106_ (
  .A(x[1]),
  .ZN(_030_)
);

NAND2_X2 _107_ (
  .A1(_029_),
  .A2(_030_),
  .ZN(_031_)
);

NAND2_X1 _108_ (
  .A1(x[2]),
  .A2(x[1]),
  .ZN(_032_)
);

NAND2_X4 _109_ (
  .A1(_031_),
  .A2(_032_),
  .ZN(_033_)
);

BUF_X4 _110_ (
  .A(y[1]),
  .Z(_034_)
);

INV_X2 _111_ (
  .A(_034_),
  .ZN(_035_)
);

AOI21_X1 _112_ (
  .A(_028_),
  .B1(_033_),
  .B2(_035_),
  .ZN(_036_)
);

INV_X1 _113_ (
  .A(x[0]),
  .ZN(_037_)
);

NAND2_X4 _114_ (
  .A1(_037_),
  .A2(_029_),
  .ZN(_038_)
);

NAND2_X1 _115_ (
  .A1(x[0]),
  .A2(x[2]),
  .ZN(_039_)
);

NAND2_X4 _116_ (
  .A1(_038_),
  .A2(_039_),
  .ZN(_040_)
);

OAI21_X1 _117_ (
  .A(_036_),
  .B1(_035_),
  .B2(_040_),
  .ZN(_041_)
);

NAND2_X1 _118_ (
  .A1(_030_),
  .A2(x[2]),
  .ZN(_042_)
);

NAND2_X2 _119_ (
  .A1(_029_),
  .A2(x[1]),
  .ZN(_043_)
);

NAND2_X4 _120_ (
  .A1(_042_),
  .A2(_043_),
  .ZN(_044_)
);

AOI21_X1 _121_ (
  .A(_027_),
  .B1(_044_),
  .B2(_034_),
  .ZN(_045_)
);

NAND2_X1 _122_ (
  .A1(_040_),
  .A2(_035_),
  .ZN(_046_)
);

NAND2_X1 _123_ (
  .A1(_045_),
  .A2(_046_),
  .ZN(_047_)
);

BUF_X1 _124_ (
  .A(ena),
  .Z(_048_)
);

BUF_X2 _125_ (
  .A(_048_),
  .Z(_049_)
);

NAND3_X1 _126_ (
  .A1(_041_),
  .A2(_047_),
  .A3(_049_),
  .ZN(_050_)
);

INV_X1 _127_ (
  .A(_048_),
  .ZN(_051_)
);

NAND2_X1 _128_ (
  .A1(_051_),
  .A2(\coef[21] ),
  .ZN(_052_)
);

NAND2_X1 _129_ (
  .A1(_050_),
  .A2(_052_),
  .ZN(_000_)
);

BUF_X2 _130_ (
  .A(y[0]),
  .Z(_053_)
);

INV_X1 _131_ (
  .A(_053_),
  .ZN(_054_)
);

NAND2_X2 _132_ (
  .A1(_040_),
  .A2(_054_),
  .ZN(_055_)
);

NAND3_X1 _133_ (
  .A1(_038_),
  .A2(_053_),
  .A3(_039_),
  .ZN(_056_)
);

NAND2_X1 _134_ (
  .A1(_055_),
  .A2(_056_),
  .ZN(_057_)
);

MUX2_X1 _135_ (
  .A(\coef[22] ),
  .B(_057_),
  .S(_048_),
  .Z(_001_)
);

NAND2_X1 _136_ (
  .A1(_033_),
  .A2(_054_),
  .ZN(_058_)
);

NAND3_X1 _137_ (
  .A1(_058_),
  .A2(_056_),
  .A3(_034_),
  .ZN(_059_)
);

NAND2_X1 _138_ (
  .A1(_059_),
  .A2(_036_),
  .ZN(_060_)
);

NAND3_X1 _139_ (
  .A1(_031_),
  .A2(_053_),
  .A3(_032_),
  .ZN(_061_)
);

NAND3_X1 _140_ (
  .A1(_055_),
  .A2(_061_),
  .A3(_035_),
  .ZN(_062_)
);

NAND2_X1 _141_ (
  .A1(_062_),
  .A2(_045_),
  .ZN(_063_)
);

NAND2_X1 _142_ (
  .A1(_060_),
  .A2(_063_),
  .ZN(_064_)
);

NAND2_X1 _143_ (
  .A1(_064_),
  .A2(_049_),
  .ZN(_065_)
);

NAND2_X1 _144_ (
  .A1(_051_),
  .A2(\coef[23] ),
  .ZN(_066_)
);

NAND2_X1 _145_ (
  .A1(_065_),
  .A2(_066_),
  .ZN(_002_)
);

NOR2_X1 _146_ (
  .A1(_049_),
  .A2(\coef[24] ),
  .ZN(_067_)
);

NAND2_X1 _147_ (
  .A1(_027_),
  .A2(_034_),
  .ZN(_068_)
);

NOR2_X1 _148_ (
  .A1(_027_),
  .A2(_034_),
  .ZN(_069_)
);

OAI21_X1 _149_ (
  .A(_068_),
  .B1(_069_),
  .B2(_053_),
  .ZN(_070_)
);

XNOR2_X1 _150_ (
  .A(_070_),
  .B(_040_),
  .ZN(_071_)
);

AOI21_X1 _151_ (
  .A(_067_),
  .B1(_071_),
  .B2(_049_),
  .ZN(_003_)
);

NAND2_X1 _152_ (
  .A1(_033_),
  .A2(_035_),
  .ZN(_072_)
);

NOR2_X1 _153_ (
  .A1(_044_),
  .A2(_028_),
  .ZN(_073_)
);

OAI21_X1 _154_ (
  .A(_072_),
  .B1(_073_),
  .B2(_069_),
  .ZN(_074_)
);

NOR2_X1 _155_ (
  .A1(_035_),
  .A2(_027_),
  .ZN(_075_)
);

NAND3_X1 _156_ (
  .A1(_058_),
  .A2(_056_),
  .A3(_075_),
  .ZN(_076_)
);

NAND2_X1 _157_ (
  .A1(_074_),
  .A2(_076_),
  .ZN(_077_)
);

NOR2_X1 _158_ (
  .A1(_028_),
  .A2(_034_),
  .ZN(_078_)
);

NAND3_X1 _159_ (
  .A1(_055_),
  .A2(_061_),
  .A3(_078_),
  .ZN(_079_)
);

NAND2_X1 _160_ (
  .A1(_079_),
  .A2(_048_),
  .ZN(_080_)
);

NOR2_X1 _161_ (
  .A1(_077_),
  .A2(_080_),
  .ZN(_081_)
);

NOR2_X1 _162_ (
  .A1(_049_),
  .A2(\coef[25] ),
  .ZN(_082_)
);

NOR2_X2 _163_ (
  .A1(_081_),
  .A2(_082_),
  .ZN(_004_)
);

OAI21_X1 _164_ (
  .A(_040_),
  .B1(_053_),
  .B2(_034_),
  .ZN(_083_)
);

NAND3_X1 _165_ (
  .A1(_033_),
  .A2(_054_),
  .A3(_035_),
  .ZN(_084_)
);

NAND3_X1 _166_ (
  .A1(_083_),
  .A2(_084_),
  .A3(_028_),
  .ZN(_085_)
);

NAND2_X1 _167_ (
  .A1(_053_),
  .A2(_034_),
  .ZN(_086_)
);

OR2_X1 _168_ (
  .A1(_033_),
  .A2(_086_),
  .ZN(_087_)
);

NAND3_X1 _169_ (
  .A1(_038_),
  .A2(_039_),
  .A3(_086_),
  .ZN(_088_)
);

NAND3_X1 _170_ (
  .A1(_087_),
  .A2(_027_),
  .A3(_088_),
  .ZN(_089_)
);

NAND2_X1 _171_ (
  .A1(_085_),
  .A2(_089_),
  .ZN(_090_)
);

NAND2_X1 _172_ (
  .A1(_090_),
  .A2(_049_),
  .ZN(_091_)
);

NAND2_X1 _173_ (
  .A1(_051_),
  .A2(\coef[26] ),
  .ZN(_092_)
);

NAND2_X1 _174_ (
  .A1(_091_),
  .A2(_092_),
  .ZN(_005_)
);

NAND2_X1 _175_ (
  .A1(_051_),
  .A2(\coef[27] ),
  .ZN(_010_)
);

NOR2_X1 _176_ (
  .A1(_078_),
  .A2(_075_),
  .ZN(_011_)
);

NAND3_X1 _177_ (
  .A1(_058_),
  .A2(_061_),
  .A3(_011_),
  .ZN(_012_)
);

NAND2_X1 _178_ (
  .A1(_012_),
  .A2(_049_),
  .ZN(_013_)
);

AOI21_X1 _179_ (
  .A(_011_),
  .B1(_055_),
  .B2(_056_),
  .ZN(_014_)
);

OAI21_X1 _180_ (
  .A(_010_),
  .B1(_013_),
  .B2(_014_),
  .ZN(_006_)
);

NAND2_X1 _181_ (
  .A1(_044_),
  .A2(_034_),
  .ZN(_015_)
);

NAND2_X1 _182_ (
  .A1(_072_),
  .A2(_015_),
  .ZN(_016_)
);

MUX2_X1 _183_ (
  .A(\coef[28] ),
  .B(_016_),
  .S(_049_),
  .Z(_007_)
);

NAND3_X1 _184_ (
  .A1(_044_),
  .A2(_054_),
  .A3(_035_),
  .ZN(_017_)
);

NAND3_X1 _185_ (
  .A1(_083_),
  .A2(_017_),
  .A3(_027_),
  .ZN(_018_)
);

OR2_X2 _186_ (
  .A1(_044_),
  .A2(_086_),
  .ZN(_019_)
);

NAND3_X1 _187_ (
  .A1(_019_),
  .A2(_028_),
  .A3(_088_),
  .ZN(_020_)
);

NAND2_X1 _188_ (
  .A1(_018_),
  .A2(_020_),
  .ZN(_021_)
);

NAND2_X1 _189_ (
  .A1(_021_),
  .A2(_049_),
  .ZN(_022_)
);

NAND2_X1 _190_ (
  .A1(_051_),
  .A2(\coef[15] ),
  .ZN(_023_)
);

NAND2_X1 _191_ (
  .A1(_022_),
  .A2(_023_),
  .ZN(_008_)
);

NOR2_X1 _192_ (
  .A1(_049_),
  .A2(\coef[30] ),
  .ZN(_024_)
);

NOR2_X1 _193_ (
  .A1(_073_),
  .A2(_051_),
  .ZN(_025_)
);

NAND2_X1 _194_ (
  .A1(_044_),
  .A2(_028_),
  .ZN(_026_)
);

AOI21_X1 _195_ (
  .A(_024_),
  .B1(_025_),
  .B2(_026_),
  .ZN(_009_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_102_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_101_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_100_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[24] ),
  .QN(_099_)
);

DFF_X1 \coef[25]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[25] ),
  .QN(_098_)
);

DFF_X1 \coef[26]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[26] ),
  .QN(_097_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[27] ),
  .QN(_096_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_095_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_094_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\coef[30] ),
  .QN(_093_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[30] , \coef[30] , \coef[15] , \coef[28] , \coef[27] , \coef[26] , \coef[25] , \coef[24] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$f5bb6813249a03e2893277297591ec050ac518dc\dctu

module \$paramod\div_su\z_width=s32'00000000000000000000000000011000 (input clk, input ena,
 input [23:0] z, input [11:0] d, output [12:0] q, output [11:0] s, output div0, output ovf);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _048_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _394_;
wire _395_;
wire _396_;
wire _397_;
wire _398_;
wire _399_;
wire _400_;
wire _401_;
wire _402_;
wire _403_;
wire _404_;
wire _405_;
wire _406_;
wire _407_;
wire _408_;
wire _409_;
wire _410_;
wire _411_;
wire _412_;
wire _413_;
wire _414_;
wire _415_;
wire _429_;
wire _431_;
wire _432_;
wire _433_;
wire _434_;
wire _435_;
wire _436_;
wire _437_;
wire _438_;
wire _439_;
wire _440_;
wire _441_;
wire _442_;
wire _443_;
wire _444_;
wire _445_;
wire _446_;
wire _447_;
wire _448_;
wire _449_;
wire _450_;
wire _451_;
wire _452_;
wire _453_;
wire _454_;
wire _455_;
wire _456_;
wire _457_;
wire _458_;
wire _459_;
wire _460_;
wire _461_;
wire _462_;
wire _463_;
wire _464_;
wire _465_;
wire _466_;
wire _467_;
wire _468_;
wire _469_;
wire _470_;
wire _471_;
wire _472_;
wire _473_;
wire _474_;
wire _475_;
wire _476_;
wire _477_;
wire _482_;
wire _483_;
wire _484_;
wire _485_;
wire _486_;
wire _487_;
wire _488_;
wire _489_;
wire \id[0] ;
wire \id[10] ;
wire \id[11] ;
wire \id[1] ;
wire \id[2] ;
wire \id[3] ;
wire \id[4] ;
wire \id[5] ;
wire \id[6] ;
wire \id[7] ;
wire \id[8] ;
wire \id[9] ;
wire idiv0;
wire iovf;
wire \iq[0] ;
wire \iq[10] ;
wire \iq[11] ;
wire \iq[1] ;
wire \iq[2] ;
wire \iq[3] ;
wire \iq[4] ;
wire \iq[5] ;
wire \iq[6] ;
wire \iq[7] ;
wire \iq[8] ;
wire \iq[9] ;
wire \is[0] ;
wire \is[10] ;
wire \is[11] ;
wire \is[1] ;
wire \is[2] ;
wire \is[3] ;
wire \is[4] ;
wire \is[5] ;
wire \is[6] ;
wire \is[7] ;
wire \is[8] ;
wire \is[9] ;
wire \iz[0] ;
wire \iz[10] ;
wire \iz[11] ;
wire \iz[12] ;
wire \iz[13] ;
wire \iz[14] ;
wire \iz[15] ;
wire \iz[16] ;
wire \iz[17] ;
wire \iz[18] ;
wire \iz[19] ;
wire \iz[1] ;
wire \iz[20] ;
wire \iz[21] ;
wire \iz[22] ;
wire \iz[23] ;
wire \iz[2] ;
wire \iz[3] ;
wire \iz[4] ;
wire \iz[5] ;
wire \iz[6] ;
wire \iz[7] ;
wire \iz[8] ;
wire \iz[9] ;
wire \spipe[0] ;
wire \spipe[10] ;
wire \spipe[11] ;
wire \spipe[12] ;
wire \spipe[13] ;
wire \spipe[1] ;
wire \spipe[2] ;
wire \spipe[3] ;
wire \spipe[4] ;
wire \spipe[5] ;
wire \spipe[6] ;
wire \spipe[7] ;
wire \spipe[8] ;
wire \spipe[9] ;

INV_X2 _490_ (
  .A(z[0]),
  .ZN(_486_)
);

INV_X1 _492_ (
  .A(\iq[0] ),
  .ZN(_482_)
);

INV_X1 _494_ (
  .A(\iq[1] ),
  .ZN(_483_)
);

INV_X2 _495_ (
  .A(z[1]),
  .ZN(_487_)
);

BUF_X1 _496_ (
  .A(ena),
  .Z(_077_)
);

INV_X1 _497_ (
  .A(_077_),
  .ZN(_078_)
);

BUF_X2 _498_ (
  .A(_078_),
  .Z(_079_)
);

NAND2_X1 _499_ (
  .A1(_079_),
  .A2(\iz[0] ),
  .ZN(_080_)
);

BUF_X2 _500_ (
  .A(_078_),
  .Z(_081_)
);

OAI21_X1 _501_ (
  .A(_080_),
  .B1(_486_),
  .B2(_081_),
  .ZN(_000_)
);

BUF_X4 _502_ (
  .A(z[23]),
  .Z(_082_)
);

INV_X4 _503_ (
  .A(_082_),
  .ZN(_083_)
);

AOI21_X1 _504_ (
  .A(_078_),
  .B1(_487_),
  .B2(_083_),
  .ZN(_084_)
);

OAI21_X1 _505_ (
  .A(_084_),
  .B1(_083_),
  .B2(_489_),
  .ZN(_085_)
);

BUF_X4 _506_ (
  .A(_077_),
  .Z(_086_)
);

BUF_X2 _507_ (
  .A(_086_),
  .Z(_087_)
);

INV_X1 _508_ (
  .A(\iz[1] ),
  .ZN(_088_)
);

OAI21_X1 _509_ (
  .A(_085_),
  .B1(_087_),
  .B2(_088_),
  .ZN(_001_)
);

BUF_X2 _510_ (
  .A(_086_),
  .Z(_089_)
);

NOR2_X1 _511_ (
  .A1(_089_),
  .A2(\iz[2] ),
  .ZN(_090_)
);

NOR2_X1 _512_ (
  .A1(_083_),
  .A2(_488_),
  .ZN(_091_)
);

XNOR2_X1 _513_ (
  .A(_091_),
  .B(z[2]),
  .ZN(_092_)
);

AOI21_X1 _514_ (
  .A(_090_),
  .B1(_092_),
  .B2(_087_),
  .ZN(_002_)
);

BUF_X2 _515_ (
  .A(_086_),
  .Z(_093_)
);

NOR2_X1 _516_ (
  .A1(_093_),
  .A2(\iz[3] ),
  .ZN(_094_)
);

INV_X2 _517_ (
  .A(z[2]),
  .ZN(_095_)
);

NAND3_X4 _518_ (
  .A1(_487_),
  .A2(_095_),
  .A3(_486_),
  .ZN(_096_)
);

BUF_X4 _519_ (
  .A(_082_),
  .Z(_097_)
);

NAND2_X1 _520_ (
  .A1(_096_),
  .A2(_097_),
  .ZN(_098_)
);

INV_X2 _521_ (
  .A(z[3]),
  .ZN(_099_)
);

XNOR2_X1 _522_ (
  .A(_098_),
  .B(_099_),
  .ZN(_100_)
);

BUF_X1 _523_ (
  .A(_086_),
  .Z(_101_)
);

AOI21_X1 _524_ (
  .A(_094_),
  .B1(_100_),
  .B2(_101_),
  .ZN(_003_)
);

BUF_X2 _525_ (
  .A(_086_),
  .Z(_102_)
);

NOR2_X1 _526_ (
  .A1(_102_),
  .A2(\iz[4] ),
  .ZN(_103_)
);

NAND3_X2 _527_ (
  .A1(_095_),
  .A2(_099_),
  .A3(_488_),
  .ZN(_104_)
);

NAND2_X2 _528_ (
  .A1(_104_),
  .A2(_082_),
  .ZN(_105_)
);

INV_X1 _529_ (
  .A(z[4]),
  .ZN(_106_)
);

XNOR2_X1 _530_ (
  .A(_105_),
  .B(_106_),
  .ZN(_107_)
);

AOI21_X1 _531_ (
  .A(_103_),
  .B1(_107_),
  .B2(_101_),
  .ZN(_004_)
);

NOR2_X1 _532_ (
  .A1(_102_),
  .A2(\iz[5] ),
  .ZN(_108_)
);

NOR2_X2 _533_ (
  .A1(z[3]),
  .A2(z[4]),
  .ZN(_109_)
);

INV_X1 _534_ (
  .A(_109_),
  .ZN(_110_)
);

NOR2_X2 _535_ (
  .A1(_096_),
  .A2(_110_),
  .ZN(_111_)
);

NOR2_X1 _536_ (
  .A1(_111_),
  .A2(_083_),
  .ZN(_112_)
);

XNOR2_X1 _537_ (
  .A(_112_),
  .B(z[5]),
  .ZN(_113_)
);

AOI21_X1 _538_ (
  .A(_108_),
  .B1(_113_),
  .B2(_101_),
  .ZN(_005_)
);

NOR2_X1 _539_ (
  .A1(_102_),
  .A2(\iz[6] ),
  .ZN(_114_)
);

NOR2_X2 _540_ (
  .A1(z[4]),
  .A2(z[5]),
  .ZN(_115_)
);

INV_X1 _541_ (
  .A(_115_),
  .ZN(_116_)
);

NOR2_X2 _542_ (
  .A1(_104_),
  .A2(_116_),
  .ZN(_117_)
);

NOR2_X1 _543_ (
  .A1(_117_),
  .A2(_083_),
  .ZN(_118_)
);

XNOR2_X1 _544_ (
  .A(_118_),
  .B(z[6]),
  .ZN(_119_)
);

AOI21_X1 _545_ (
  .A(_114_),
  .B1(_119_),
  .B2(_101_),
  .ZN(_006_)
);

NOR2_X1 _546_ (
  .A1(_093_),
  .A2(\iz[7] ),
  .ZN(_120_)
);

NOR2_X2 _547_ (
  .A1(z[5]),
  .A2(z[6]),
  .ZN(_121_)
);

NAND2_X2 _548_ (
  .A1(_109_),
  .A2(_121_),
  .ZN(_122_)
);

NOR2_X4 _549_ (
  .A1(_122_),
  .A2(_096_),
  .ZN(_123_)
);

NOR2_X1 _550_ (
  .A1(_123_),
  .A2(_083_),
  .ZN(_124_)
);

XNOR2_X1 _551_ (
  .A(_124_),
  .B(z[7]),
  .ZN(_125_)
);

AOI21_X1 _552_ (
  .A(_120_),
  .B1(_125_),
  .B2(_101_),
  .ZN(_007_)
);

NOR2_X1 _553_ (
  .A1(_102_),
  .A2(\iz[8] ),
  .ZN(_126_)
);

NOR2_X2 _554_ (
  .A1(z[6]),
  .A2(z[7]),
  .ZN(_127_)
);

NAND2_X1 _555_ (
  .A1(_115_),
  .A2(_127_),
  .ZN(_128_)
);

NAND2_X2 _556_ (
  .A1(_128_),
  .A2(_082_),
  .ZN(_129_)
);

NAND2_X4 _557_ (
  .A1(_129_),
  .A2(_105_),
  .ZN(_130_)
);

XNOR2_X1 _558_ (
  .A(_130_),
  .B(z[8]),
  .ZN(_131_)
);

BUF_X2 _559_ (
  .A(_086_),
  .Z(_132_)
);

AOI21_X1 _560_ (
  .A(_126_),
  .B1(_131_),
  .B2(_132_),
  .ZN(_008_)
);

CLKBUF_X3 _561_ (
  .A(_086_),
  .Z(_133_)
);

NOR2_X1 _562_ (
  .A1(_133_),
  .A2(\iz[9] ),
  .ZN(_134_)
);

NOR2_X2 _563_ (
  .A1(z[7]),
  .A2(z[8]),
  .ZN(_135_)
);

NAND2_X1 _564_ (
  .A1(_123_),
  .A2(_135_),
  .ZN(_136_)
);

NAND2_X2 _565_ (
  .A1(_136_),
  .A2(_082_),
  .ZN(_137_)
);

INV_X1 _566_ (
  .A(z[9]),
  .ZN(_138_)
);

XNOR2_X2 _567_ (
  .A(_137_),
  .B(_138_),
  .ZN(_139_)
);

AOI21_X2 _568_ (
  .A(_134_),
  .B1(_139_),
  .B2(_132_),
  .ZN(_009_)
);

NOR2_X1 _569_ (
  .A1(_093_),
  .A2(\iz[10] ),
  .ZN(_140_)
);

NOR2_X2 _570_ (
  .A1(z[8]),
  .A2(z[9]),
  .ZN(_141_)
);

NOR2_X1 _571_ (
  .A1(_141_),
  .A2(_083_),
  .ZN(_142_)
);

INV_X1 _572_ (
  .A(_142_),
  .ZN(_143_)
);

NAND3_X2 _573_ (
  .A1(_129_),
  .A2(_105_),
  .A3(_143_),
  .ZN(_144_)
);

XNOR2_X1 _574_ (
  .A(_144_),
  .B(z[10]),
  .ZN(_145_)
);

AOI21_X1 _575_ (
  .A(_140_),
  .B1(_145_),
  .B2(_132_),
  .ZN(_010_)
);

NOR2_X1 _576_ (
  .A1(_089_),
  .A2(\iz[11] ),
  .ZN(_146_)
);

NOR2_X2 _577_ (
  .A1(z[9]),
  .A2(z[10]),
  .ZN(_147_)
);

AND2_X1 _578_ (
  .A1(_135_),
  .A2(_147_),
  .ZN(_148_)
);

NAND2_X1 _579_ (
  .A1(_123_),
  .A2(_148_),
  .ZN(_149_)
);

NAND2_X2 _580_ (
  .A1(_149_),
  .A2(_082_),
  .ZN(_150_)
);

INV_X1 _581_ (
  .A(z[11]),
  .ZN(_151_)
);

XNOR2_X2 _582_ (
  .A(_150_),
  .B(_151_),
  .ZN(_152_)
);

AOI21_X2 _583_ (
  .A(_146_),
  .B1(_152_),
  .B2(_132_),
  .ZN(_011_)
);

NOR2_X1 _584_ (
  .A1(_089_),
  .A2(\iz[12] ),
  .ZN(_153_)
);

NOR2_X2 _585_ (
  .A1(z[10]),
  .A2(z[11]),
  .ZN(_154_)
);

NAND2_X1 _586_ (
  .A1(_141_),
  .A2(_154_),
  .ZN(_155_)
);

NAND2_X1 _587_ (
  .A1(_155_),
  .A2(_082_),
  .ZN(_156_)
);

INV_X1 _588_ (
  .A(_156_),
  .ZN(_157_)
);

NOR2_X4 _589_ (
  .A1(_130_),
  .A2(_157_),
  .ZN(_158_)
);

INV_X1 _590_ (
  .A(z[12]),
  .ZN(_159_)
);

XNOR2_X2 _591_ (
  .A(_158_),
  .B(_159_),
  .ZN(_160_)
);

AOI21_X2 _592_ (
  .A(_153_),
  .B1(_160_),
  .B2(_101_),
  .ZN(_012_)
);

NOR2_X1 _593_ (
  .A1(_133_),
  .A2(\iz[13] ),
  .ZN(_161_)
);

NAND2_X1 _594_ (
  .A1(_121_),
  .A2(_135_),
  .ZN(_162_)
);

NOR2_X2 _595_ (
  .A1(z[11]),
  .A2(z[12]),
  .ZN(_163_)
);

NAND2_X2 _596_ (
  .A1(_147_),
  .A2(_163_),
  .ZN(_164_)
);

NOR2_X2 _597_ (
  .A1(_162_),
  .A2(_164_),
  .ZN(_165_)
);

NAND2_X1 _598_ (
  .A1(_165_),
  .A2(_111_),
  .ZN(_166_)
);

NAND2_X2 _599_ (
  .A1(_166_),
  .A2(_082_),
  .ZN(_167_)
);

INV_X1 _600_ (
  .A(z[13]),
  .ZN(_168_)
);

XNOR2_X2 _601_ (
  .A(_167_),
  .B(_168_),
  .ZN(_169_)
);

AOI21_X2 _602_ (
  .A(_161_),
  .B1(_169_),
  .B2(_087_),
  .ZN(_013_)
);

NOR2_X1 _603_ (
  .A1(_089_),
  .A2(\iz[14] ),
  .ZN(_170_)
);

NOR2_X2 _604_ (
  .A1(z[12]),
  .A2(z[13]),
  .ZN(_171_)
);

NAND2_X1 _605_ (
  .A1(_127_),
  .A2(_171_),
  .ZN(_172_)
);

NOR2_X1 _606_ (
  .A1(_155_),
  .A2(_172_),
  .ZN(_173_)
);

NAND2_X1 _607_ (
  .A1(_173_),
  .A2(_117_),
  .ZN(_174_)
);

NAND2_X2 _608_ (
  .A1(_174_),
  .A2(_097_),
  .ZN(_175_)
);

INV_X1 _609_ (
  .A(z[14]),
  .ZN(_176_)
);

XNOR2_X2 _610_ (
  .A(_175_),
  .B(_176_),
  .ZN(_177_)
);

AOI21_X2 _611_ (
  .A(_170_),
  .B1(_177_),
  .B2(_132_),
  .ZN(_014_)
);

NOR2_X1 _612_ (
  .A1(_089_),
  .A2(\iz[15] ),
  .ZN(_178_)
);

NAND2_X1 _613_ (
  .A1(_135_),
  .A2(_147_),
  .ZN(_179_)
);

NOR2_X2 _614_ (
  .A1(z[13]),
  .A2(z[14]),
  .ZN(_180_)
);

NAND2_X1 _615_ (
  .A1(_163_),
  .A2(_180_),
  .ZN(_181_)
);

NOR2_X1 _616_ (
  .A1(_179_),
  .A2(_181_),
  .ZN(_182_)
);

NAND2_X1 _617_ (
  .A1(_182_),
  .A2(_123_),
  .ZN(_183_)
);

NAND2_X2 _618_ (
  .A1(_183_),
  .A2(_097_),
  .ZN(_184_)
);

INV_X1 _619_ (
  .A(z[15]),
  .ZN(_185_)
);

XNOR2_X2 _620_ (
  .A(_184_),
  .B(_185_),
  .ZN(_186_)
);

AOI21_X2 _621_ (
  .A(_178_),
  .B1(_186_),
  .B2(_087_),
  .ZN(_015_)
);

NOR2_X1 _622_ (
  .A1(z[14]),
  .A2(z[15]),
  .ZN(_187_)
);

NAND2_X1 _623_ (
  .A1(_171_),
  .A2(_187_),
  .ZN(_188_)
);

NAND2_X1 _624_ (
  .A1(_188_),
  .A2(_097_),
  .ZN(_189_)
);

NAND2_X1 _625_ (
  .A1(_158_),
  .A2(_189_),
  .ZN(_190_)
);

NAND2_X1 _626_ (
  .A1(_190_),
  .A2(z[16]),
  .ZN(_191_)
);

INV_X1 _627_ (
  .A(z[16]),
  .ZN(_192_)
);

NAND3_X1 _628_ (
  .A1(_158_),
  .A2(_192_),
  .A3(_189_),
  .ZN(_193_)
);

NAND3_X1 _629_ (
  .A1(_191_),
  .A2(_193_),
  .A3(_133_),
  .ZN(_194_)
);

NAND2_X1 _630_ (
  .A1(_081_),
  .A2(\iz[16] ),
  .ZN(_195_)
);

NAND2_X1 _631_ (
  .A1(_194_),
  .A2(_195_),
  .ZN(_016_)
);

NOR2_X1 _632_ (
  .A1(z[15]),
  .A2(z[16]),
  .ZN(_196_)
);

NAND2_X1 _633_ (
  .A1(_180_),
  .A2(_196_),
  .ZN(_197_)
);

OAI21_X1 _634_ (
  .A(_097_),
  .B1(_164_),
  .B2(_197_),
  .ZN(_198_)
);

NAND2_X1 _635_ (
  .A1(_137_),
  .A2(_198_),
  .ZN(_199_)
);

NAND2_X1 _636_ (
  .A1(_199_),
  .A2(z[17]),
  .ZN(_200_)
);

INV_X1 _637_ (
  .A(z[17]),
  .ZN(_201_)
);

NAND3_X1 _638_ (
  .A1(_137_),
  .A2(_201_),
  .A3(_198_),
  .ZN(_202_)
);

NAND3_X1 _639_ (
  .A1(_200_),
  .A2(_202_),
  .A3(_133_),
  .ZN(_203_)
);

NAND2_X1 _640_ (
  .A1(_081_),
  .A2(\iz[17] ),
  .ZN(_204_)
);

NAND2_X1 _641_ (
  .A1(_203_),
  .A2(_204_),
  .ZN(_017_)
);

INV_X1 _642_ (
  .A(_144_),
  .ZN(_205_)
);

NAND2_X1 _643_ (
  .A1(_154_),
  .A2(_171_),
  .ZN(_206_)
);

NOR2_X1 _644_ (
  .A1(z[16]),
  .A2(z[17]),
  .ZN(_207_)
);

NAND2_X1 _645_ (
  .A1(_187_),
  .A2(_207_),
  .ZN(_208_)
);

OAI21_X1 _646_ (
  .A(_097_),
  .B1(_206_),
  .B2(_208_),
  .ZN(_209_)
);

NAND2_X1 _647_ (
  .A1(_205_),
  .A2(_209_),
  .ZN(_210_)
);

NAND2_X1 _648_ (
  .A1(_210_),
  .A2(z[18]),
  .ZN(_211_)
);

INV_X1 _649_ (
  .A(z[18]),
  .ZN(_212_)
);

NAND3_X1 _650_ (
  .A1(_205_),
  .A2(_212_),
  .A3(_209_),
  .ZN(_213_)
);

NAND3_X1 _651_ (
  .A1(_211_),
  .A2(_213_),
  .A3(_133_),
  .ZN(_214_)
);

NAND2_X1 _652_ (
  .A1(_081_),
  .A2(\iz[18] ),
  .ZN(_215_)
);

NAND2_X1 _653_ (
  .A1(_214_),
  .A2(_215_),
  .ZN(_018_)
);

NOR2_X1 _654_ (
  .A1(z[17]),
  .A2(z[18]),
  .ZN(_216_)
);

NAND2_X1 _655_ (
  .A1(_196_),
  .A2(_216_),
  .ZN(_217_)
);

OAI21_X1 _656_ (
  .A(_097_),
  .B1(_181_),
  .B2(_217_),
  .ZN(_218_)
);

NAND2_X1 _657_ (
  .A1(_150_),
  .A2(_218_),
  .ZN(_219_)
);

NAND2_X1 _658_ (
  .A1(_219_),
  .A2(z[19]),
  .ZN(_220_)
);

INV_X1 _659_ (
  .A(z[19]),
  .ZN(_221_)
);

NAND3_X1 _660_ (
  .A1(_150_),
  .A2(_221_),
  .A3(_218_),
  .ZN(_222_)
);

NAND3_X1 _661_ (
  .A1(_220_),
  .A2(_222_),
  .A3(_133_),
  .ZN(_223_)
);

NAND2_X1 _662_ (
  .A1(_079_),
  .A2(\iz[19] ),
  .ZN(_224_)
);

NAND2_X1 _663_ (
  .A1(_223_),
  .A2(_224_),
  .ZN(_019_)
);

NOR2_X1 _664_ (
  .A1(z[18]),
  .A2(z[19]),
  .ZN(_225_)
);

NAND2_X1 _665_ (
  .A1(_207_),
  .A2(_225_),
  .ZN(_226_)
);

OAI21_X1 _666_ (
  .A(_097_),
  .B1(_188_),
  .B2(_226_),
  .ZN(_227_)
);

NAND2_X1 _667_ (
  .A1(_158_),
  .A2(_227_),
  .ZN(_228_)
);

NAND2_X1 _668_ (
  .A1(_228_),
  .A2(z[20]),
  .ZN(_229_)
);

INV_X1 _669_ (
  .A(z[20]),
  .ZN(_230_)
);

NAND3_X1 _670_ (
  .A1(_158_),
  .A2(_230_),
  .A3(_227_),
  .ZN(_231_)
);

CLKBUF_X3 _671_ (
  .A(_086_),
  .Z(_232_)
);

NAND3_X1 _672_ (
  .A1(_229_),
  .A2(_231_),
  .A3(_232_),
  .ZN(_233_)
);

NAND2_X1 _673_ (
  .A1(_081_),
  .A2(\iz[20] ),
  .ZN(_234_)
);

NAND2_X1 _674_ (
  .A1(_233_),
  .A2(_234_),
  .ZN(_020_)
);

NOR2_X1 _675_ (
  .A1(z[19]),
  .A2(z[20]),
  .ZN(_235_)
);

NAND2_X1 _676_ (
  .A1(_180_),
  .A2(_235_),
  .ZN(_236_)
);

OAI21_X1 _677_ (
  .A(_097_),
  .B1(_217_),
  .B2(_236_),
  .ZN(_237_)
);

NAND2_X1 _678_ (
  .A1(_167_),
  .A2(_237_),
  .ZN(_238_)
);

NAND2_X1 _679_ (
  .A1(_238_),
  .A2(z[21]),
  .ZN(_239_)
);

INV_X1 _680_ (
  .A(z[21]),
  .ZN(_240_)
);

NAND3_X1 _681_ (
  .A1(_167_),
  .A2(_240_),
  .A3(_237_),
  .ZN(_241_)
);

NAND3_X1 _682_ (
  .A1(_239_),
  .A2(_241_),
  .A3(_232_),
  .ZN(_242_)
);

NAND2_X1 _683_ (
  .A1(_079_),
  .A2(\iz[21] ),
  .ZN(_243_)
);

NAND2_X1 _684_ (
  .A1(_242_),
  .A2(_243_),
  .ZN(_021_)
);

NOR2_X1 _685_ (
  .A1(z[20]),
  .A2(z[21]),
  .ZN(_244_)
);

NAND2_X1 _686_ (
  .A1(_225_),
  .A2(_244_),
  .ZN(_245_)
);

OAI21_X1 _687_ (
  .A(_097_),
  .B1(_208_),
  .B2(_245_),
  .ZN(_246_)
);

NAND2_X1 _688_ (
  .A1(_175_),
  .A2(_246_),
  .ZN(_247_)
);

NAND2_X1 _689_ (
  .A1(_247_),
  .A2(z[22]),
  .ZN(_248_)
);

INV_X1 _690_ (
  .A(z[22]),
  .ZN(_249_)
);

NAND3_X1 _691_ (
  .A1(_175_),
  .A2(_249_),
  .A3(_246_),
  .ZN(_250_)
);

NAND3_X1 _692_ (
  .A1(_248_),
  .A2(_250_),
  .A3(_232_),
  .ZN(_251_)
);

NAND2_X1 _693_ (
  .A1(_079_),
  .A2(\iz[22] ),
  .ZN(_252_)
);

NAND2_X1 _694_ (
  .A1(_251_),
  .A2(_252_),
  .ZN(_022_)
);

NAND2_X1 _695_ (
  .A1(_078_),
  .A2(q[0]),
  .ZN(_253_)
);

OAI21_X1 _696_ (
  .A(_253_),
  .B1(_482_),
  .B2(_081_),
  .ZN(_023_)
);

CLKBUF_X2 _697_ (
  .A(\spipe[13] ),
  .Z(_254_)
);

INV_X2 _698_ (
  .A(_254_),
  .ZN(_255_)
);

AOI21_X1 _699_ (
  .A(_078_),
  .B1(_483_),
  .B2(_255_),
  .ZN(_256_)
);

OAI21_X1 _700_ (
  .A(_256_),
  .B1(_255_),
  .B2(_485_),
  .ZN(_257_)
);

INV_X1 _701_ (
  .A(q[1]),
  .ZN(_258_)
);

OAI21_X1 _702_ (
  .A(_257_),
  .B1(_087_),
  .B2(_258_),
  .ZN(_024_)
);

NOR2_X1 _703_ (
  .A1(_093_),
  .A2(q[2]),
  .ZN(_259_)
);

INV_X1 _704_ (
  .A(_484_),
  .ZN(_260_)
);

BUF_X4 _705_ (
  .A(_254_),
  .Z(_261_)
);

NAND2_X1 _706_ (
  .A1(_260_),
  .A2(_261_),
  .ZN(_262_)
);

INV_X1 _707_ (
  .A(\iq[2] ),
  .ZN(_263_)
);

XNOR2_X1 _708_ (
  .A(_262_),
  .B(_263_),
  .ZN(_264_)
);

AOI21_X1 _709_ (
  .A(_259_),
  .B1(_264_),
  .B2(_087_),
  .ZN(_025_)
);

NOR2_X1 _710_ (
  .A1(_089_),
  .A2(q[3]),
  .ZN(_265_)
);

NAND3_X1 _711_ (
  .A1(_263_),
  .A2(_483_),
  .A3(_482_),
  .ZN(_266_)
);

NAND2_X1 _712_ (
  .A1(_266_),
  .A2(_261_),
  .ZN(_267_)
);

INV_X1 _713_ (
  .A(\iq[3] ),
  .ZN(_268_)
);

XNOR2_X1 _714_ (
  .A(_267_),
  .B(_268_),
  .ZN(_269_)
);

AOI21_X1 _715_ (
  .A(_265_),
  .B1(_269_),
  .B2(_087_),
  .ZN(_026_)
);

NOR2_X1 _716_ (
  .A1(_089_),
  .A2(q[4]),
  .ZN(_270_)
);

NOR2_X1 _717_ (
  .A1(_260_),
  .A2(\iq[2] ),
  .ZN(_271_)
);

AOI21_X1 _718_ (
  .A(_255_),
  .B1(_271_),
  .B2(_268_),
  .ZN(_272_)
);

XNOR2_X1 _719_ (
  .A(_272_),
  .B(\iq[4] ),
  .ZN(_273_)
);

AOI21_X1 _720_ (
  .A(_270_),
  .B1(_273_),
  .B2(_132_),
  .ZN(_027_)
);

NOR2_X1 _721_ (
  .A1(_089_),
  .A2(q[5]),
  .ZN(_274_)
);

INV_X1 _722_ (
  .A(\iq[4] ),
  .ZN(_275_)
);

NAND2_X1 _723_ (
  .A1(_275_),
  .A2(_268_),
  .ZN(_276_)
);

OAI21_X1 _724_ (
  .A(_261_),
  .B1(_266_),
  .B2(_276_),
  .ZN(_277_)
);

INV_X1 _725_ (
  .A(\iq[5] ),
  .ZN(_278_)
);

XNOR2_X1 _726_ (
  .A(_277_),
  .B(_278_),
  .ZN(_279_)
);

AOI21_X1 _727_ (
  .A(_274_),
  .B1(_279_),
  .B2(_132_),
  .ZN(_028_)
);

NOR2_X1 _728_ (
  .A1(_089_),
  .A2(q[6]),
  .ZN(_280_)
);

NOR2_X2 _729_ (
  .A1(\iq[4] ),
  .A2(\iq[3] ),
  .ZN(_281_)
);

NAND3_X1 _730_ (
  .A1(_271_),
  .A2(_281_),
  .A3(_278_),
  .ZN(_282_)
);

NAND2_X1 _731_ (
  .A1(_282_),
  .A2(_261_),
  .ZN(_283_)
);

INV_X1 _732_ (
  .A(\iq[6] ),
  .ZN(_284_)
);

XNOR2_X1 _733_ (
  .A(_283_),
  .B(_284_),
  .ZN(_285_)
);

AOI21_X1 _734_ (
  .A(_280_),
  .B1(_285_),
  .B2(_132_),
  .ZN(_029_)
);

NOR2_X1 _735_ (
  .A1(_089_),
  .A2(q[7]),
  .ZN(_286_)
);

NAND3_X1 _736_ (
  .A1(_281_),
  .A2(_284_),
  .A3(_278_),
  .ZN(_287_)
);

NOR2_X2 _737_ (
  .A1(_287_),
  .A2(_266_),
  .ZN(_288_)
);

NOR2_X1 _738_ (
  .A1(_288_),
  .A2(_255_),
  .ZN(_289_)
);

BUF_X1 _739_ (
  .A(\iq[7] ),
  .Z(_290_)
);

XNOR2_X1 _740_ (
  .A(_289_),
  .B(_290_),
  .ZN(_291_)
);

AOI21_X1 _741_ (
  .A(_286_),
  .B1(_291_),
  .B2(_101_),
  .ZN(_030_)
);

INV_X1 _742_ (
  .A(_287_),
  .ZN(_292_)
);

NOR3_X1 _743_ (
  .A1(_260_),
  .A2(_290_),
  .A3(\iq[2] ),
  .ZN(_293_)
);

NAND2_X1 _744_ (
  .A1(_292_),
  .A2(_293_),
  .ZN(_294_)
);

BUF_X2 _745_ (
  .A(_254_),
  .Z(_295_)
);

NAND2_X1 _746_ (
  .A1(_294_),
  .A2(_295_),
  .ZN(_296_)
);

INV_X1 _747_ (
  .A(\iq[8] ),
  .ZN(_297_)
);

NAND2_X1 _748_ (
  .A1(_296_),
  .A2(_297_),
  .ZN(_298_)
);

NAND3_X1 _749_ (
  .A1(_294_),
  .A2(\iq[8] ),
  .A3(_295_),
  .ZN(_299_)
);

NAND3_X1 _750_ (
  .A1(_298_),
  .A2(_299_),
  .A3(_133_),
  .ZN(_300_)
);

INV_X1 _751_ (
  .A(q[8]),
  .ZN(_301_)
);

OAI21_X1 _752_ (
  .A(_300_),
  .B1(_087_),
  .B2(_301_),
  .ZN(_031_)
);

NOR2_X1 _753_ (
  .A1(\iq[8] ),
  .A2(_290_),
  .ZN(_302_)
);

NAND2_X1 _754_ (
  .A1(_288_),
  .A2(_302_),
  .ZN(_303_)
);

NAND2_X1 _755_ (
  .A1(_303_),
  .A2(_295_),
  .ZN(_304_)
);

INV_X1 _756_ (
  .A(\iq[9] ),
  .ZN(_305_)
);

NAND2_X1 _757_ (
  .A1(_304_),
  .A2(_305_),
  .ZN(_306_)
);

NAND3_X1 _758_ (
  .A1(_303_),
  .A2(\iq[9] ),
  .A3(_295_),
  .ZN(_307_)
);

NAND3_X1 _759_ (
  .A1(_306_),
  .A2(_307_),
  .A3(_133_),
  .ZN(_308_)
);

NAND2_X1 _760_ (
  .A1(_079_),
  .A2(q[9]),
  .ZN(_309_)
);

NAND2_X1 _761_ (
  .A1(_308_),
  .A2(_309_),
  .ZN(_032_)
);

NAND2_X1 _762_ (
  .A1(_305_),
  .A2(_297_),
  .ZN(_310_)
);

INV_X1 _763_ (
  .A(_310_),
  .ZN(_311_)
);

NAND3_X1 _764_ (
  .A1(_292_),
  .A2(_293_),
  .A3(_311_),
  .ZN(_312_)
);

NAND2_X1 _765_ (
  .A1(_312_),
  .A2(_295_),
  .ZN(_313_)
);

INV_X1 _766_ (
  .A(\iq[10] ),
  .ZN(_314_)
);

NAND2_X1 _767_ (
  .A1(_313_),
  .A2(_314_),
  .ZN(_315_)
);

NAND3_X1 _768_ (
  .A1(_312_),
  .A2(\iq[10] ),
  .A3(_295_),
  .ZN(_316_)
);

NAND3_X1 _769_ (
  .A1(_315_),
  .A2(_316_),
  .A3(_232_),
  .ZN(_317_)
);

NAND2_X1 _770_ (
  .A1(_079_),
  .A2(q[10]),
  .ZN(_318_)
);

NAND2_X1 _771_ (
  .A1(_317_),
  .A2(_318_),
  .ZN(_033_)
);

NOR3_X1 _772_ (
  .A1(_310_),
  .A2(\iq[10] ),
  .A3(_290_),
  .ZN(_319_)
);

NAND2_X1 _773_ (
  .A1(_288_),
  .A2(_319_),
  .ZN(_320_)
);

NAND2_X1 _774_ (
  .A1(_320_),
  .A2(_295_),
  .ZN(_321_)
);

INV_X1 _775_ (
  .A(\iq[11] ),
  .ZN(_322_)
);

NAND2_X1 _776_ (
  .A1(_321_),
  .A2(_322_),
  .ZN(_323_)
);

NAND3_X1 _777_ (
  .A1(_320_),
  .A2(\iq[11] ),
  .A3(_295_),
  .ZN(_324_)
);

NAND3_X1 _778_ (
  .A1(_323_),
  .A2(_324_),
  .A3(_232_),
  .ZN(_325_)
);

NAND2_X1 _779_ (
  .A1(_081_),
  .A2(q[11]),
  .ZN(_326_)
);

NAND2_X1 _780_ (
  .A1(_325_),
  .A2(_326_),
  .ZN(_034_)
);

BUF_X2 _781_ (
  .A(_077_),
  .Z(_327_)
);

MUX2_X1 _782_ (
  .A(\id[0] ),
  .B(d[0]),
  .S(_327_),
  .Z(_035_)
);

MUX2_X1 _783_ (
  .A(\id[1] ),
  .B(d[1]),
  .S(_086_),
  .Z(_036_)
);

BUF_X2 _784_ (
  .A(_086_),
  .Z(_328_)
);

MUX2_X1 _785_ (
  .A(\id[2] ),
  .B(d[2]),
  .S(_328_),
  .Z(_037_)
);

MUX2_X1 _786_ (
  .A(\id[3] ),
  .B(d[3]),
  .S(_328_),
  .Z(_038_)
);

MUX2_X1 _787_ (
  .A(\id[4] ),
  .B(d[4]),
  .S(_328_),
  .Z(_039_)
);

MUX2_X1 _788_ (
  .A(\id[5] ),
  .B(d[5]),
  .S(_328_),
  .Z(_040_)
);

MUX2_X1 _789_ (
  .A(\id[6] ),
  .B(d[6]),
  .S(_328_),
  .Z(_041_)
);

MUX2_X1 _790_ (
  .A(\id[7] ),
  .B(d[7]),
  .S(_328_),
  .Z(_042_)
);

MUX2_X1 _791_ (
  .A(\id[8] ),
  .B(d[8]),
  .S(_328_),
  .Z(_043_)
);

MUX2_X1 _792_ (
  .A(\id[9] ),
  .B(d[9]),
  .S(_328_),
  .Z(_044_)
);

MUX2_X1 _793_ (
  .A(\id[10] ),
  .B(d[10]),
  .S(_093_),
  .Z(_045_)
);

MUX2_X1 _794_ (
  .A(\id[11] ),
  .B(d[11]),
  .S(_093_),
  .Z(_046_)
);

NOR2_X1 _796_ (
  .A1(_102_),
  .A2(q[12]),
  .ZN(_329_)
);

NAND3_X1 _797_ (
  .A1(_311_),
  .A2(_322_),
  .A3(_314_),
  .ZN(_330_)
);

AOI21_X1 _798_ (
  .A(_078_),
  .B1(_330_),
  .B2(_295_),
  .ZN(_331_)
);

AOI21_X1 _799_ (
  .A(_329_),
  .B1(_331_),
  .B2(_296_),
  .ZN(_048_)
);

NAND2_X1 _875_ (
  .A1(_079_),
  .A2(\iz[23] ),
  .ZN(_394_)
);

NAND2_X1 _876_ (
  .A1(_082_),
  .A2(_077_),
  .ZN(_395_)
);

NOR3_X1 _877_ (
  .A1(_217_),
  .A2(z[21]),
  .A3(_395_),
  .ZN(_396_)
);

NAND3_X1 _878_ (
  .A1(_396_),
  .A2(_249_),
  .A3(_235_),
  .ZN(_397_)
);

OAI21_X1 _879_ (
  .A(_394_),
  .B1(_397_),
  .B2(_183_),
  .ZN(_062_)
);

INV_X1 _880_ (
  .A(\spipe[0] ),
  .ZN(_398_)
);

OAI21_X1 _881_ (
  .A(_395_),
  .B1(_087_),
  .B2(_398_),
  .ZN(_063_)
);

NAND2_X1 _882_ (
  .A1(_079_),
  .A2(\spipe[1] ),
  .ZN(_399_)
);

OAI21_X1 _883_ (
  .A(_399_),
  .B1(_081_),
  .B2(_398_),
  .ZN(_064_)
);

MUX2_X1 _884_ (
  .A(\spipe[2] ),
  .B(\spipe[1] ),
  .S(_327_),
  .Z(_065_)
);

MUX2_X1 _885_ (
  .A(\spipe[3] ),
  .B(\spipe[2] ),
  .S(_327_),
  .Z(_066_)
);

MUX2_X1 _886_ (
  .A(\spipe[4] ),
  .B(\spipe[3] ),
  .S(_327_),
  .Z(_067_)
);

MUX2_X1 _887_ (
  .A(\spipe[5] ),
  .B(\spipe[4] ),
  .S(_327_),
  .Z(_068_)
);

MUX2_X1 _888_ (
  .A(\spipe[6] ),
  .B(\spipe[5] ),
  .S(_327_),
  .Z(_069_)
);

MUX2_X1 _889_ (
  .A(\spipe[7] ),
  .B(\spipe[6] ),
  .S(_327_),
  .Z(_070_)
);

MUX2_X1 _890_ (
  .A(\spipe[8] ),
  .B(\spipe[7] ),
  .S(_327_),
  .Z(_071_)
);

MUX2_X1 _891_ (
  .A(\spipe[9] ),
  .B(\spipe[8] ),
  .S(_327_),
  .Z(_072_)
);

MUX2_X1 _892_ (
  .A(\spipe[10] ),
  .B(\spipe[9] ),
  .S(_327_),
  .Z(_073_)
);

MUX2_X1 _893_ (
  .A(\spipe[11] ),
  .B(\spipe[10] ),
  .S(_093_),
  .Z(_074_)
);

MUX2_X1 _894_ (
  .A(\spipe[12] ),
  .B(\spipe[11] ),
  .S(_328_),
  .Z(_075_)
);

NAND2_X1 _895_ (
  .A1(_232_),
  .A2(\spipe[12] ),
  .ZN(_400_)
);

OAI21_X1 _896_ (
  .A(_400_),
  .B1(_255_),
  .B2(_232_),
  .ZN(_076_)
);

HA_X1 _898_ (
  .A(_482_),
  .B(_483_),
  .CO(_484_),
  .S(_485_)
);

HA_X1 _899_ (
  .A(_486_),
  .B(_487_),
  .CO(_488_),
  .S(_489_)
);

\$paramod$ee2aa8736952ca7eee7f4751cab786a479da4583\div_uu  divider (
  .clk(clk),
  .ena(ena),
  .z({\iz[23] , \iz[22] , \iz[21] , \iz[20] , \iz[19] , \iz[18] , \iz[17] , \iz[16] , \iz[15] , \iz[14] , \iz[13] , \iz[12] , \iz[11] , \iz[10] , \iz[9] , \iz[8] , \iz[7] , \iz[6] , \iz[5] , \iz[4] , \iz[3] , \iz[2] , \iz[1] , \iz[0] }),
  .d({\id[11] , \id[10] , \id[9] , \id[8] , \id[7] , \id[6] , \id[5] , \id[4] , \id[3] , \id[2] , \id[1] , \id[0] }),
  .q({\iq[11] , \iq[10] , \iq[9] , \iq[8] , \iq[7] , \iq[6] , \iq[5] , \iq[4] , \iq[3] , \iq[2] , \iq[1] , \iq[0] }),
  .s({\is[11] , \is[10] , \is[9] , \is[8] , \is[7] , \is[6] , \is[5] , \is[4] , \is[3] , \is[2] , \is[1] , \is[0] }),
  .div0(idiv0),
  .ovf(iovf)
);

DFF_X1 \id[0]$_DFFE_PP_  (
  .D(_035_),
  .CK(clk),
  .Q(\id[0] ),
  .QN(_442_)
);

DFF_X1 \id[10]$_DFFE_PP_  (
  .D(_045_),
  .CK(clk),
  .Q(\id[10] ),
  .QN(_432_)
);

DFF_X1 \id[11]$_DFFE_PP_  (
  .D(_046_),
  .CK(clk),
  .Q(\id[11] ),
  .QN(_431_)
);

DFF_X1 \id[1]$_DFFE_PP_  (
  .D(_036_),
  .CK(clk),
  .Q(\id[1] ),
  .QN(_441_)
);

DFF_X1 \id[2]$_DFFE_PP_  (
  .D(_037_),
  .CK(clk),
  .Q(\id[2] ),
  .QN(_440_)
);

DFF_X1 \id[3]$_DFFE_PP_  (
  .D(_038_),
  .CK(clk),
  .Q(\id[3] ),
  .QN(_439_)
);

DFF_X1 \id[4]$_DFFE_PP_  (
  .D(_039_),
  .CK(clk),
  .Q(\id[4] ),
  .QN(_438_)
);

DFF_X1 \id[5]$_DFFE_PP_  (
  .D(_040_),
  .CK(clk),
  .Q(\id[5] ),
  .QN(_437_)
);

DFF_X1 \id[6]$_DFFE_PP_  (
  .D(_041_),
  .CK(clk),
  .Q(\id[6] ),
  .QN(_436_)
);

DFF_X1 \id[7]$_DFFE_PP_  (
  .D(_042_),
  .CK(clk),
  .Q(\id[7] ),
  .QN(_435_)
);

DFF_X1 \id[8]$_DFFE_PP_  (
  .D(_043_),
  .CK(clk),
  .Q(\id[8] ),
  .QN(_434_)
);

DFF_X1 \id[9]$_DFFE_PP_  (
  .D(_044_),
  .CK(clk),
  .Q(\id[9] ),
  .QN(_433_)
);

DFF_X1 \iz[0]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\iz[0] ),
  .QN(_477_)
);

DFF_X1 \iz[10]$_DFFE_PP_  (
  .D(_010_),
  .CK(clk),
  .Q(\iz[10] ),
  .QN(_467_)
);

DFF_X1 \iz[11]$_DFFE_PP_  (
  .D(_011_),
  .CK(clk),
  .Q(\iz[11] ),
  .QN(_466_)
);

DFF_X1 \iz[12]$_DFFE_PP_  (
  .D(_012_),
  .CK(clk),
  .Q(\iz[12] ),
  .QN(_465_)
);

DFF_X1 \iz[13]$_DFFE_PP_  (
  .D(_013_),
  .CK(clk),
  .Q(\iz[13] ),
  .QN(_464_)
);

DFF_X1 \iz[14]$_DFFE_PP_  (
  .D(_014_),
  .CK(clk),
  .Q(\iz[14] ),
  .QN(_463_)
);

DFF_X1 \iz[15]$_DFFE_PP_  (
  .D(_015_),
  .CK(clk),
  .Q(\iz[15] ),
  .QN(_462_)
);

DFF_X1 \iz[16]$_DFFE_PP_  (
  .D(_016_),
  .CK(clk),
  .Q(\iz[16] ),
  .QN(_461_)
);

DFF_X1 \iz[17]$_DFFE_PP_  (
  .D(_017_),
  .CK(clk),
  .Q(\iz[17] ),
  .QN(_460_)
);

DFF_X1 \iz[18]$_DFFE_PP_  (
  .D(_018_),
  .CK(clk),
  .Q(\iz[18] ),
  .QN(_459_)
);

DFF_X1 \iz[19]$_DFFE_PP_  (
  .D(_019_),
  .CK(clk),
  .Q(\iz[19] ),
  .QN(_458_)
);

DFF_X1 \iz[1]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\iz[1] ),
  .QN(_476_)
);

DFF_X1 \iz[20]$_DFFE_PP_  (
  .D(_020_),
  .CK(clk),
  .Q(\iz[20] ),
  .QN(_457_)
);

DFF_X1 \iz[21]$_DFFE_PP_  (
  .D(_021_),
  .CK(clk),
  .Q(\iz[21] ),
  .QN(_456_)
);

DFF_X1 \iz[22]$_DFFE_PP_  (
  .D(_022_),
  .CK(clk),
  .Q(\iz[22] ),
  .QN(_455_)
);

DFF_X1 \iz[23]$_SDFFCE_PN0P_  (
  .D(_062_),
  .CK(clk),
  .Q(\iz[23] ),
  .QN(_415_)
);

DFF_X1 \iz[2]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\iz[2] ),
  .QN(_475_)
);

DFF_X1 \iz[3]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\iz[3] ),
  .QN(_474_)
);

DFF_X1 \iz[4]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\iz[4] ),
  .QN(_473_)
);

DFF_X1 \iz[5]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\iz[5] ),
  .QN(_472_)
);

DFF_X1 \iz[6]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\iz[6] ),
  .QN(_471_)
);

DFF_X1 \iz[7]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\iz[7] ),
  .QN(_470_)
);

DFF_X1 \iz[8]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(\iz[8] ),
  .QN(_469_)
);

DFF_X1 \iz[9]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(\iz[9] ),
  .QN(_468_)
);

DFF_X1 \q[0]$_DFFE_PP_  (
  .D(_023_),
  .CK(clk),
  .Q(q[0]),
  .QN(_454_)
);

DFF_X1 \q[10]$_DFFE_PP_  (
  .D(_033_),
  .CK(clk),
  .Q(q[10]),
  .QN(_444_)
);

DFF_X1 \q[11]$_DFFE_PP_  (
  .D(_034_),
  .CK(clk),
  .Q(q[11]),
  .QN(_443_)
);

DFF_X1 \q[12]$_SDFFCE_PN0P_  (
  .D(_048_),
  .CK(clk),
  .Q(q[12]),
  .QN(_429_)
);

DFF_X1 \q[1]$_DFFE_PP_  (
  .D(_024_),
  .CK(clk),
  .Q(q[1]),
  .QN(_453_)
);

DFF_X1 \q[2]$_DFFE_PP_  (
  .D(_025_),
  .CK(clk),
  .Q(q[2]),
  .QN(_452_)
);

DFF_X1 \q[3]$_DFFE_PP_  (
  .D(_026_),
  .CK(clk),
  .Q(q[3]),
  .QN(_451_)
);

DFF_X1 \q[4]$_DFFE_PP_  (
  .D(_027_),
  .CK(clk),
  .Q(q[4]),
  .QN(_450_)
);

DFF_X1 \q[5]$_DFFE_PP_  (
  .D(_028_),
  .CK(clk),
  .Q(q[5]),
  .QN(_449_)
);

DFF_X1 \q[6]$_DFFE_PP_  (
  .D(_029_),
  .CK(clk),
  .Q(q[6]),
  .QN(_448_)
);

DFF_X1 \q[7]$_DFFE_PP_  (
  .D(_030_),
  .CK(clk),
  .Q(q[7]),
  .QN(_447_)
);

DFF_X1 \q[8]$_DFFE_PP_  (
  .D(_031_),
  .CK(clk),
  .Q(q[8]),
  .QN(_446_)
);

DFF_X1 \q[9]$_DFFE_PP_  (
  .D(_032_),
  .CK(clk),
  .Q(q[9]),
  .QN(_445_)
);

DFF_X1 \spipe[0]$_DFFE_PP_  (
  .D(_063_),
  .CK(clk),
  .Q(\spipe[0] ),
  .QN(_414_)
);

DFF_X1 \spipe[10]$_DFFE_PP_  (
  .D(_073_),
  .CK(clk),
  .Q(\spipe[10] ),
  .QN(_404_)
);

DFF_X1 \spipe[11]$_DFFE_PP_  (
  .D(_074_),
  .CK(clk),
  .Q(\spipe[11] ),
  .QN(_403_)
);

DFF_X1 \spipe[12]$_DFFE_PP_  (
  .D(_075_),
  .CK(clk),
  .Q(\spipe[12] ),
  .QN(_402_)
);

DFF_X1 \spipe[13]$_DFFE_PP_  (
  .D(_076_),
  .CK(clk),
  .Q(\spipe[13] ),
  .QN(_401_)
);

DFF_X1 \spipe[1]$_DFFE_PP_  (
  .D(_064_),
  .CK(clk),
  .Q(\spipe[1] ),
  .QN(_413_)
);

DFF_X1 \spipe[2]$_DFFE_PP_  (
  .D(_065_),
  .CK(clk),
  .Q(\spipe[2] ),
  .QN(_412_)
);

DFF_X1 \spipe[3]$_DFFE_PP_  (
  .D(_066_),
  .CK(clk),
  .Q(\spipe[3] ),
  .QN(_411_)
);

DFF_X1 \spipe[4]$_DFFE_PP_  (
  .D(_067_),
  .CK(clk),
  .Q(\spipe[4] ),
  .QN(_410_)
);

DFF_X1 \spipe[5]$_DFFE_PP_  (
  .D(_068_),
  .CK(clk),
  .Q(\spipe[5] ),
  .QN(_409_)
);

DFF_X1 \spipe[6]$_DFFE_PP_  (
  .D(_069_),
  .CK(clk),
  .Q(\spipe[6] ),
  .QN(_408_)
);

DFF_X1 \spipe[7]$_DFFE_PP_  (
  .D(_070_),
  .CK(clk),
  .Q(\spipe[7] ),
  .QN(_407_)
);

DFF_X1 \spipe[8]$_DFFE_PP_  (
  .D(_071_),
  .CK(clk),
  .Q(\spipe[8] ),
  .QN(_406_)
);

DFF_X1 \spipe[9]$_DFFE_PP_  (
  .D(_072_),
  .CK(clk),
  .Q(\spipe[9] ),
  .QN(_405_)
);
endmodule //$paramod\div_su\z_width=s32'00000000000000000000000000011000

module \$paramod$f878842d6bc0ac80c3f795bb76ef86af701fb0a2\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _069_ (
  .A(x[0]),
  .ZN(_051_)
);

INV_X1 _070_ (
  .A(x[1]),
  .ZN(_052_)
);

BUF_X4 _071_ (
  .A(ena),
  .Z(_008_)
);

INV_X4 _072_ (
  .A(_008_),
  .ZN(_009_)
);

NAND2_X1 _073_ (
  .A1(_009_),
  .A2(\coef[21] ),
  .ZN(_010_)
);

OAI21_X1 _074_ (
  .A(_010_),
  .B1(x[1]),
  .B2(_009_),
  .ZN(_000_)
);

NAND2_X1 _075_ (
  .A1(_009_),
  .A2(\coef[22] ),
  .ZN(_011_)
);

BUF_X4 _076_ (
  .A(x[2]),
  .Z(_012_)
);

NAND2_X1 _077_ (
  .A1(_012_),
  .A2(_053_),
  .ZN(_013_)
);

NAND2_X1 _078_ (
  .A1(_013_),
  .A2(_008_),
  .ZN(_014_)
);

NOR2_X1 _079_ (
  .A1(_067_),
  .A2(_012_),
  .ZN(_015_)
);

OAI21_X1 _080_ (
  .A(_011_),
  .B1(_014_),
  .B2(_015_),
  .ZN(_001_)
);

INV_X1 _081_ (
  .A(_059_),
  .ZN(_016_)
);

NAND2_X1 _082_ (
  .A1(_016_),
  .A2(_012_),
  .ZN(_017_)
);

INV_X4 _083_ (
  .A(_012_),
  .ZN(_018_)
);

NAND2_X1 _084_ (
  .A1(_018_),
  .A2(_061_),
  .ZN(_019_)
);

NAND3_X1 _085_ (
  .A1(_017_),
  .A2(_019_),
  .A3(_008_),
  .ZN(_020_)
);

NAND2_X1 _086_ (
  .A1(_009_),
  .A2(\coef[23] ),
  .ZN(_021_)
);

NAND2_X1 _087_ (
  .A1(_020_),
  .A2(_021_),
  .ZN(_002_)
);

INV_X1 _088_ (
  .A(_055_),
  .ZN(_022_)
);

NAND2_X1 _089_ (
  .A1(_022_),
  .A2(_012_),
  .ZN(_023_)
);

NAND2_X1 _090_ (
  .A1(_018_),
  .A2(_065_),
  .ZN(_024_)
);

NAND3_X1 _091_ (
  .A1(_023_),
  .A2(_024_),
  .A3(_008_),
  .ZN(_025_)
);

NAND2_X1 _092_ (
  .A1(_009_),
  .A2(\coef[14] ),
  .ZN(_026_)
);

NAND2_X1 _093_ (
  .A1(_025_),
  .A2(_026_),
  .ZN(_003_)
);

NAND2_X1 _094_ (
  .A1(_009_),
  .A2(\coef[13] ),
  .ZN(_027_)
);

OAI21_X1 _095_ (
  .A(_027_),
  .B1(_018_),
  .B2(_009_),
  .ZN(_004_)
);

INV_X1 _096_ (
  .A(_054_),
  .ZN(_028_)
);

NAND2_X1 _097_ (
  .A1(_018_),
  .A2(_028_),
  .ZN(_029_)
);

NAND2_X1 _098_ (
  .A1(_012_),
  .A2(_054_),
  .ZN(_030_)
);

NAND3_X1 _099_ (
  .A1(_029_),
  .A2(_008_),
  .A3(_030_),
  .ZN(_031_)
);

NAND2_X1 _100_ (
  .A1(_009_),
  .A2(\coef[28] ),
  .ZN(_032_)
);

NAND2_X1 _101_ (
  .A1(_031_),
  .A2(_032_),
  .ZN(_005_)
);

INV_X1 _102_ (
  .A(_063_),
  .ZN(_033_)
);

NAND2_X1 _103_ (
  .A1(_033_),
  .A2(_012_),
  .ZN(_034_)
);

NAND2_X1 _104_ (
  .A1(_018_),
  .A2(_057_),
  .ZN(_035_)
);

NAND3_X1 _105_ (
  .A1(_034_),
  .A2(_035_),
  .A3(_008_),
  .ZN(_036_)
);

NAND2_X1 _106_ (
  .A1(_009_),
  .A2(\coef[15] ),
  .ZN(_037_)
);

NAND2_X1 _107_ (
  .A1(_036_),
  .A2(_037_),
  .ZN(_006_)
);

INV_X1 _108_ (
  .A(_067_),
  .ZN(_038_)
);

NAND2_X1 _109_ (
  .A1(_038_),
  .A2(_012_),
  .ZN(_039_)
);

NAND2_X1 _110_ (
  .A1(_018_),
  .A2(_053_),
  .ZN(_040_)
);

NAND3_X1 _111_ (
  .A1(_039_),
  .A2(_040_),
  .A3(_008_),
  .ZN(_041_)
);

NAND2_X1 _112_ (
  .A1(_009_),
  .A2(\coef[12] ),
  .ZN(_042_)
);

NAND2_X1 _113_ (
  .A1(_041_),
  .A2(_042_),
  .ZN(_007_)
);

HA_X1 _114_ (
  .A(_051_),
  .B(_052_),
  .CO(_053_),
  .S(_054_)
);

HA_X1 _115_ (
  .A(_051_),
  .B(_052_),
  .CO(_055_),
  .S(_056_)
);

HA_X1 _116_ (
  .A(_051_),
  .B(x[1]),
  .CO(_057_),
  .S(_058_)
);

HA_X1 _117_ (
  .A(_051_),
  .B(x[1]),
  .CO(_059_),
  .S(_060_)
);

HA_X1 _118_ (
  .A(x[0]),
  .B(_052_),
  .CO(_061_),
  .S(_062_)
);

HA_X1 _119_ (
  .A(x[0]),
  .B(_052_),
  .CO(_063_),
  .S(_064_)
);

HA_X1 _120_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_065_),
  .S(_066_)
);

HA_X1 _121_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_067_),
  .S(_068_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_050_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_049_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_048_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_047_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_046_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_045_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_044_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_043_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$f878842d6bc0ac80c3f795bb76ef86af701fb0a2\dctu

module \$paramod$fa41e4d02884503da5d6c381e868b8c261424a31\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire \coef[10] ;
wire \coef[11] ;
wire \coef[13] ;
wire \coef[15] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

NOR2_X1 _34_ (
  .A1(\coef[11] ),
  .A2(ena),
  .ZN(_04_)
);

INV_X1 _35_ (
  .A(ena),
  .ZN(_05_)
);

INV_X1 _36_ (
  .A(x[1]),
  .ZN(_06_)
);

INV_X1 _37_ (
  .A(x[0]),
  .ZN(_07_)
);

NAND2_X2 _38_ (
  .A1(_06_),
  .A2(_07_),
  .ZN(_08_)
);

NAND2_X1 _39_ (
  .A1(x[1]),
  .A2(x[0]),
  .ZN(_09_)
);

NAND2_X4 _40_ (
  .A1(_08_),
  .A2(_09_),
  .ZN(_10_)
);

INV_X1 _41_ (
  .A(y[1]),
  .ZN(_11_)
);

INV_X2 _42_ (
  .A(y[2]),
  .ZN(_12_)
);

NAND2_X4 _43_ (
  .A1(_11_),
  .A2(_12_),
  .ZN(_13_)
);

NAND2_X1 _44_ (
  .A1(y[1]),
  .A2(y[2]),
  .ZN(_14_)
);

NAND2_X4 _45_ (
  .A1(_13_),
  .A2(_14_),
  .ZN(_15_)
);

AOI21_X4 _46_ (
  .A(_05_),
  .B1(_10_),
  .B2(_15_),
  .ZN(_16_)
);

OR2_X4 _47_ (
  .A1(_15_),
  .A2(_10_),
  .ZN(_17_)
);

AOI21_X4 _48_ (
  .A(_04_),
  .B1(_16_),
  .B2(_17_),
  .ZN(_00_)
);

XNOR2_X2 _49_ (
  .A(_12_),
  .B(y[0]),
  .ZN(_18_)
);

INV_X2 _50_ (
  .A(_10_),
  .ZN(_19_)
);

NAND2_X2 _51_ (
  .A1(_18_),
  .A2(_19_),
  .ZN(_20_)
);

XNOR2_X1 _52_ (
  .A(y[2]),
  .B(y[0]),
  .ZN(_21_)
);

NAND2_X1 _53_ (
  .A1(_21_),
  .A2(_10_),
  .ZN(_22_)
);

NAND3_X1 _54_ (
  .A1(_20_),
  .A2(_22_),
  .A3(ena),
  .ZN(_23_)
);

NAND2_X1 _55_ (
  .A1(_05_),
  .A2(\coef[13] ),
  .ZN(_24_)
);

NAND2_X1 _56_ (
  .A1(_23_),
  .A2(_24_),
  .ZN(_01_)
);

NAND2_X1 _57_ (
  .A1(_20_),
  .A2(_22_),
  .ZN(_25_)
);

NAND2_X1 _58_ (
  .A1(_25_),
  .A2(ena),
  .ZN(_26_)
);

NAND2_X1 _59_ (
  .A1(_05_),
  .A2(\coef[10] ),
  .ZN(_27_)
);

NAND2_X1 _60_ (
  .A1(_26_),
  .A2(_27_),
  .ZN(_02_)
);

NAND2_X4 _61_ (
  .A1(_16_),
  .A2(_17_),
  .ZN(_28_)
);

NAND2_X1 _62_ (
  .A1(_05_),
  .A2(\coef[15] ),
  .ZN(_29_)
);

NAND2_X2 _63_ (
  .A1(_28_),
  .A2(_29_),
  .ZN(_03_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\coef[11] ),
  .QN(_33_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_01_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_32_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_02_),
  .CK(clk),
  .Q(\coef[10] ),
  .QN(_31_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_03_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_30_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[15] , \coef[15] , \coef[10] , \coef[13] , \coef[10] , \coef[15] , \coef[15] , \coef[11] , \coef[10] , \coef[11] , \coef[15] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$fa41e4d02884503da5d6c381e868b8c261424a31\dctu

module \$paramod$1b119bd029c81aaa2221a23d15ab3b6b02f6efee\dctu (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire \coef[12] ;
wire \coef[13] ;
wire \coef[14] ;
wire \coef[15] ;
wire \coef[21] ;
wire \coef[22] ;
wire \coef[23] ;
wire \coef[28] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;

INV_X1 _116_ (
  .A(x[0]),
  .ZN(_098_)
);

INV_X1 _117_ (
  .A(x[1]),
  .ZN(_099_)
);

BUF_X4 _118_ (
  .A(x[2]),
  .Z(_032_)
);

NAND2_X1 _119_ (
  .A1(_101_),
  .A2(_032_),
  .ZN(_033_)
);

INV_X1 _120_ (
  .A(_033_),
  .ZN(_034_)
);

BUF_X16 _121_ (
  .A(_032_),
  .Z(_035_)
);

NOR2_X4 _122_ (
  .A1(_101_),
  .A2(_035_),
  .ZN(_036_)
);

NOR2_X2 _123_ (
  .A1(_034_),
  .A2(_036_),
  .ZN(_037_)
);

XNOR2_X2 _124_ (
  .A(y[0]),
  .B(y[1]),
  .ZN(_038_)
);

NAND2_X1 _125_ (
  .A1(_037_),
  .A2(_038_),
  .ZN(_039_)
);

INV_X1 _126_ (
  .A(_101_),
  .ZN(_040_)
);

INV_X4 _127_ (
  .A(_032_),
  .ZN(_041_)
);

NAND2_X1 _128_ (
  .A1(_040_),
  .A2(_041_),
  .ZN(_042_)
);

NAND2_X1 _129_ (
  .A1(_042_),
  .A2(_033_),
  .ZN(_043_)
);

INV_X1 _130_ (
  .A(y[0]),
  .ZN(_044_)
);

NAND2_X1 _131_ (
  .A1(_044_),
  .A2(y[1]),
  .ZN(_045_)
);

INV_X1 _132_ (
  .A(y[1]),
  .ZN(_046_)
);

NAND2_X1 _133_ (
  .A1(_046_),
  .A2(y[0]),
  .ZN(_047_)
);

NAND2_X2 _134_ (
  .A1(_045_),
  .A2(_047_),
  .ZN(_048_)
);

NAND2_X1 _135_ (
  .A1(_043_),
  .A2(_048_),
  .ZN(_049_)
);

BUF_X2 _136_ (
  .A(ena),
  .Z(_050_)
);

NAND3_X1 _137_ (
  .A1(_039_),
  .A2(_049_),
  .A3(_050_),
  .ZN(_051_)
);

INV_X1 _138_ (
  .A(_050_),
  .ZN(_052_)
);

NAND2_X1 _139_ (
  .A1(_052_),
  .A2(\coef[21] ),
  .ZN(_053_)
);

NAND2_X1 _140_ (
  .A1(_051_),
  .A2(_053_),
  .ZN(_000_)
);

INV_X1 _141_ (
  .A(_106_),
  .ZN(_054_)
);

NAND2_X1 _142_ (
  .A1(_041_),
  .A2(_054_),
  .ZN(_055_)
);

NAND2_X2 _143_ (
  .A1(_035_),
  .A2(_108_),
  .ZN(_056_)
);

NAND2_X1 _144_ (
  .A1(_055_),
  .A2(_056_),
  .ZN(_057_)
);

NAND2_X1 _145_ (
  .A1(_038_),
  .A2(_057_),
  .ZN(_058_)
);

NAND2_X1 _146_ (
  .A1(_041_),
  .A2(_104_),
  .ZN(_059_)
);

INV_X1 _147_ (
  .A(_110_),
  .ZN(_060_)
);

NAND2_X2 _148_ (
  .A1(_060_),
  .A2(_035_),
  .ZN(_061_)
);

NAND2_X2 _149_ (
  .A1(_059_),
  .A2(_061_),
  .ZN(_062_)
);

NAND2_X1 _150_ (
  .A1(_048_),
  .A2(_062_),
  .ZN(_063_)
);

NAND3_X1 _151_ (
  .A1(_058_),
  .A2(_063_),
  .A3(_050_),
  .ZN(_064_)
);

NAND2_X1 _152_ (
  .A1(_052_),
  .A2(\coef[22] ),
  .ZN(_065_)
);

NAND2_X1 _153_ (
  .A1(_064_),
  .A2(_065_),
  .ZN(_001_)
);

NAND2_X4 _154_ (
  .A1(_035_),
  .A2(_114_),
  .ZN(_066_)
);

INV_X2 _155_ (
  .A(_066_),
  .ZN(_067_)
);

NOR2_X2 _156_ (
  .A1(_035_),
  .A2(_100_),
  .ZN(_068_)
);

NOR2_X2 _157_ (
  .A1(_067_),
  .A2(_068_),
  .ZN(_069_)
);

NAND2_X1 _158_ (
  .A1(_069_),
  .A2(_038_),
  .ZN(_070_)
);

INV_X1 _159_ (
  .A(_102_),
  .ZN(_071_)
);

NAND2_X1 _160_ (
  .A1(_041_),
  .A2(_071_),
  .ZN(_072_)
);

NAND2_X1 _161_ (
  .A1(_035_),
  .A2(_112_),
  .ZN(_073_)
);

NAND2_X1 _162_ (
  .A1(_072_),
  .A2(_073_),
  .ZN(_074_)
);

NAND2_X1 _163_ (
  .A1(_048_),
  .A2(_074_),
  .ZN(_075_)
);

NAND3_X1 _164_ (
  .A1(_070_),
  .A2(_075_),
  .A3(_050_),
  .ZN(_076_)
);

NAND2_X1 _165_ (
  .A1(_052_),
  .A2(\coef[23] ),
  .ZN(_077_)
);

NAND2_X1 _166_ (
  .A1(_076_),
  .A2(_077_),
  .ZN(_002_)
);

NAND2_X1 _167_ (
  .A1(_038_),
  .A2(_062_),
  .ZN(_078_)
);

NAND2_X1 _168_ (
  .A1(_048_),
  .A2(_057_),
  .ZN(_079_)
);

NAND3_X1 _169_ (
  .A1(_078_),
  .A2(_079_),
  .A3(_050_),
  .ZN(_080_)
);

NAND2_X1 _170_ (
  .A1(_052_),
  .A2(\coef[14] ),
  .ZN(_081_)
);

NAND2_X1 _171_ (
  .A1(_080_),
  .A2(_081_),
  .ZN(_003_)
);

NAND2_X1 _172_ (
  .A1(_038_),
  .A2(x[0]),
  .ZN(_082_)
);

NAND2_X1 _173_ (
  .A1(_048_),
  .A2(_098_),
  .ZN(_083_)
);

NAND3_X1 _174_ (
  .A1(_082_),
  .A2(_083_),
  .A3(_050_),
  .ZN(_084_)
);

NAND2_X1 _175_ (
  .A1(_052_),
  .A2(\coef[13] ),
  .ZN(_085_)
);

NAND2_X1 _176_ (
  .A1(_084_),
  .A2(_085_),
  .ZN(_004_)
);

NAND2_X1 _177_ (
  .A1(_038_),
  .A2(x[1]),
  .ZN(_086_)
);

NAND2_X1 _178_ (
  .A1(_048_),
  .A2(_099_),
  .ZN(_087_)
);

NAND3_X1 _179_ (
  .A1(_086_),
  .A2(_087_),
  .A3(_050_),
  .ZN(_088_)
);

NAND2_X1 _180_ (
  .A1(_052_),
  .A2(\coef[28] ),
  .ZN(_089_)
);

NAND2_X1 _181_ (
  .A1(_088_),
  .A2(_089_),
  .ZN(_005_)
);

NAND2_X1 _182_ (
  .A1(_041_),
  .A2(_114_),
  .ZN(_008_)
);

INV_X1 _183_ (
  .A(_100_),
  .ZN(_009_)
);

NAND2_X4 _184_ (
  .A1(_009_),
  .A2(_035_),
  .ZN(_010_)
);

NAND2_X2 _185_ (
  .A1(_008_),
  .A2(_010_),
  .ZN(_011_)
);

INV_X1 _186_ (
  .A(_011_),
  .ZN(_012_)
);

NAND2_X1 _187_ (
  .A1(_012_),
  .A2(_038_),
  .ZN(_013_)
);

NAND2_X1 _188_ (
  .A1(_041_),
  .A2(_112_),
  .ZN(_014_)
);

NAND2_X1 _189_ (
  .A1(_071_),
  .A2(_035_),
  .ZN(_015_)
);

NAND2_X1 _190_ (
  .A1(_014_),
  .A2(_015_),
  .ZN(_016_)
);

NAND2_X1 _191_ (
  .A1(_048_),
  .A2(_016_),
  .ZN(_017_)
);

NAND3_X1 _192_ (
  .A1(_013_),
  .A2(_017_),
  .A3(_050_),
  .ZN(_018_)
);

NAND2_X1 _193_ (
  .A1(_052_),
  .A2(\coef[15] ),
  .ZN(_019_)
);

NAND2_X1 _194_ (
  .A1(_018_),
  .A2(_019_),
  .ZN(_006_)
);

NAND2_X1 _195_ (
  .A1(_041_),
  .A2(_110_),
  .ZN(_020_)
);

INV_X1 _196_ (
  .A(_104_),
  .ZN(_021_)
);

NAND2_X4 _197_ (
  .A1(_021_),
  .A2(_035_),
  .ZN(_022_)
);

NAND2_X2 _198_ (
  .A1(_020_),
  .A2(_022_),
  .ZN(_023_)
);

INV_X1 _199_ (
  .A(_023_),
  .ZN(_024_)
);

NAND2_X1 _200_ (
  .A1(_024_),
  .A2(_038_),
  .ZN(_025_)
);

NAND2_X1 _201_ (
  .A1(_041_),
  .A2(_108_),
  .ZN(_026_)
);

NAND2_X1 _202_ (
  .A1(_054_),
  .A2(_035_),
  .ZN(_027_)
);

NAND2_X1 _203_ (
  .A1(_026_),
  .A2(_027_),
  .ZN(_028_)
);

NAND2_X1 _204_ (
  .A1(_048_),
  .A2(_028_),
  .ZN(_029_)
);

NAND3_X1 _205_ (
  .A1(_025_),
  .A2(_029_),
  .A3(_050_),
  .ZN(_030_)
);

NAND2_X1 _206_ (
  .A1(_052_),
  .A2(\coef[12] ),
  .ZN(_031_)
);

NAND2_X1 _207_ (
  .A1(_030_),
  .A2(_031_),
  .ZN(_007_)
);

HA_X1 _208_ (
  .A(_098_),
  .B(_099_),
  .CO(_100_),
  .S(_101_)
);

HA_X1 _209_ (
  .A(_098_),
  .B(_099_),
  .CO(_102_),
  .S(_103_)
);

HA_X1 _210_ (
  .A(_098_),
  .B(x[1]),
  .CO(_104_),
  .S(_105_)
);

HA_X1 _211_ (
  .A(_098_),
  .B(x[1]),
  .CO(_106_),
  .S(_107_)
);

HA_X1 _212_ (
  .A(x[0]),
  .B(_099_),
  .CO(_108_),
  .S(_109_)
);

HA_X1 _213_ (
  .A(x[0]),
  .B(_099_),
  .CO(_110_),
  .S(_111_)
);

HA_X1 _214_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_112_),
  .S(_113_)
);

HA_X1 _215_ (
  .A(x[0]),
  .B(x[1]),
  .CO(_114_),
  .S(_115_)
);

DFF_X1 \coef[21]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(\coef[21] ),
  .QN(_097_)
);

DFF_X1 \coef[22]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(\coef[22] ),
  .QN(_096_)
);

DFF_X1 \coef[23]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(\coef[23] ),
  .QN(_095_)
);

DFF_X1 \coef[24]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(\coef[14] ),
  .QN(_094_)
);

DFF_X1 \coef[27]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(\coef[13] ),
  .QN(_093_)
);

DFF_X1 \coef[28]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(\coef[28] ),
  .QN(_092_)
);

DFF_X1 \coef[29]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(\coef[15] ),
  .QN(_091_)
);

DFF_X1 \coef[31]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(\coef[12] ),
  .QN(_090_)
);

\$paramod$b5a8bcf0c5a3eb6704410e66fd72520afc96ea51\dct_mac  macu (
  .clk(clk),
  .ena(ena),
  .dclr(ddgo),
  .din(ddin),
  .coef({\coef[12] , \coef[12] , \coef[15] , \coef[28] , \coef[13] , \coef[15] , \coef[12] , \coef[14] , \coef[23] , \coef[22] , \coef[21] }),
  .result({dout, \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
);
endmodule //$paramod$1b119bd029c81aaa2221a23d15ab3b6b02f6efee\dctu

module \$paramod$f79433e3440244ebaeb06fcd795abd5555024789\dctub (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout0, output [11:0] dout1,
 output [11:0] dout2, output [11:0] dout3, output [11:0] dout4, output [11:0] dout5, output [11:0] dout6,
 output [11:0] dout7);
\$paramod$8cd9bf70556f3aa976ca66d64ee3b9c1b3a94e21\dctu  dct_unit_0 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout0)
);

\$paramod$30e2d72cbb2d6c7d2f48769e891fec5593e1f756\dctu  dct_unit_1 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout1)
);

\$paramod$022e4835c44d221125856d68f8603b7186431212\dctu  dct_unit_2 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout2)
);

\$paramod$f878842d6bc0ac80c3f795bb76ef86af701fb0a2\dctu  dct_unit_3 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout3)
);

\$paramod$bd5d8b7ea001bd9da1e8d07da4940a1f4c75e6b0\dctu  dct_unit_4 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout4)
);

\$paramod$bb43d9c07810ea45f23a5f680ee116bafcd9334e\dctu  dct_unit_5 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout5)
);

\$paramod$c50cce30a10e9eb82ea37b86647b55ab680286c8\dctu  dct_unit_6 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout6)
);

\$paramod$9f831900faf0e9bfdbd9e0f8aa853df59256a109\dctu  dct_unit_7 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout7)
);
endmodule //$paramod$f79433e3440244ebaeb06fcd795abd5555024789\dctub

module jpeg_qnr(input clk, input ena, input rst, input dstrb, input [11:0] din, input [7:0] qnt_val,
 output [5:0] qnt_cnt, output [10:0] dout, output douten);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire \dep[0] ;
wire \dep[10] ;
wire \dep[11] ;
wire \dep[12] ;
wire \dep[13] ;
wire \dep[14] ;
wire \dep[1] ;
wire \dep[2] ;
wire \dep[3] ;
wire \dep[4] ;
wire \dep[5] ;
wire \dep[6] ;
wire \dep[7] ;
wire \dep[8] ;
wire \dep[9] ;
wire \iq[0] ;
wire \iq[10] ;
wire \iq[11] ;
wire \iq[12] ;
wire \iq[1] ;
wire \iq[2] ;
wire \iq[3] ;
wire \iq[4] ;
wire \iq[5] ;
wire \iq[6] ;
wire \iq[7] ;
wire \iq[8] ;
wire \iq[9] ;

BUF_X4 _294_ (
  .A(ena),
  .Z(_033_)
);

INV_X1 _295_ (
  .A(_033_),
  .ZN(_034_)
);

BUF_X2 _296_ (
  .A(_034_),
  .Z(_035_)
);

NAND2_X1 _297_ (
  .A1(_035_),
  .A2(dout[0]),
  .ZN(_036_)
);

BUF_X4 _298_ (
  .A(\iq[0] ),
  .Z(_037_)
);

NAND2_X4 _299_ (
  .A1(_037_),
  .A2(_272_),
  .ZN(_038_)
);

BUF_X2 _300_ (
  .A(_033_),
  .Z(_039_)
);

NAND2_X1 _301_ (
  .A1(_038_),
  .A2(_039_),
  .ZN(_040_)
);

BUF_X2 _302_ (
  .A(_037_),
  .Z(_041_)
);

NOR2_X1 _303_ (
  .A1(_041_),
  .A2(\iq[1] ),
  .ZN(_042_)
);

OAI21_X1 _304_ (
  .A(_036_),
  .B1(_040_),
  .B2(_042_),
  .ZN(_000_)
);

NAND2_X1 _305_ (
  .A1(_035_),
  .A2(dout[1]),
  .ZN(_043_)
);

INV_X1 _306_ (
  .A(_271_),
  .ZN(_044_)
);

NAND2_X4 _307_ (
  .A1(_038_),
  .A2(_044_),
  .ZN(_045_)
);

INV_X4 _308_ (
  .A(_045_),
  .ZN(_046_)
);

BUF_X4 _309_ (
  .A(_274_),
  .Z(_047_)
);

XNOR2_X1 _310_ (
  .A(_046_),
  .B(_047_),
  .ZN(_048_)
);

INV_X2 _311_ (
  .A(_037_),
  .ZN(_049_)
);

OAI21_X1 _312_ (
  .A(_039_),
  .B1(_048_),
  .B2(_049_),
  .ZN(_050_)
);

NOR2_X1 _313_ (
  .A1(_041_),
  .A2(\iq[2] ),
  .ZN(_051_)
);

OAI21_X1 _314_ (
  .A(_043_),
  .B1(_050_),
  .B2(_051_),
  .ZN(_001_)
);

NAND2_X1 _315_ (
  .A1(_035_),
  .A2(dout[2]),
  .ZN(_052_)
);

NAND2_X4 _316_ (
  .A1(_047_),
  .A2(_271_),
  .ZN(_053_)
);

INV_X1 _317_ (
  .A(_273_),
  .ZN(_054_)
);

NAND2_X2 _318_ (
  .A1(_053_),
  .A2(_054_),
  .ZN(_055_)
);

INV_X2 _319_ (
  .A(_055_),
  .ZN(_056_)
);

NAND2_X4 _320_ (
  .A1(_047_),
  .A2(_272_),
  .ZN(_057_)
);

INV_X4 _321_ (
  .A(_057_),
  .ZN(_058_)
);

NAND2_X2 _322_ (
  .A1(_058_),
  .A2(_037_),
  .ZN(_059_)
);

NAND2_X2 _323_ (
  .A1(_056_),
  .A2(_059_),
  .ZN(_060_)
);

INV_X1 _324_ (
  .A(_060_),
  .ZN(_061_)
);

BUF_X4 _325_ (
  .A(_276_),
  .Z(_062_)
);

XNOR2_X1 _326_ (
  .A(_061_),
  .B(_062_),
  .ZN(_063_)
);

OAI21_X1 _327_ (
  .A(_039_),
  .B1(_063_),
  .B2(_049_),
  .ZN(_064_)
);

NOR2_X1 _328_ (
  .A1(_041_),
  .A2(\iq[3] ),
  .ZN(_065_)
);

OAI21_X2 _329_ (
  .A(_052_),
  .B1(_064_),
  .B2(_065_),
  .ZN(_002_)
);

INV_X1 _330_ (
  .A(\iq[4] ),
  .ZN(_066_)
);

OAI21_X1 _331_ (
  .A(_033_),
  .B1(_066_),
  .B2(_037_),
  .ZN(_067_)
);

NAND2_X4 _332_ (
  .A1(_062_),
  .A2(_273_),
  .ZN(_068_)
);

INV_X1 _333_ (
  .A(_275_),
  .ZN(_069_)
);

NAND2_X2 _334_ (
  .A1(_068_),
  .A2(_069_),
  .ZN(_070_)
);

INV_X1 _335_ (
  .A(_070_),
  .ZN(_071_)
);

NAND2_X4 _336_ (
  .A1(_047_),
  .A2(_062_),
  .ZN(_072_)
);

OAI21_X4 _337_ (
  .A(_071_),
  .B1(_046_),
  .B2(_072_),
  .ZN(_073_)
);

BUF_X4 _338_ (
  .A(_278_),
  .Z(_074_)
);

XOR2_X2 _339_ (
  .A(_073_),
  .B(_074_),
  .Z(_075_)
);

AOI21_X2 _340_ (
  .A(_067_),
  .B1(_075_),
  .B2(_041_),
  .ZN(_076_)
);

NOR2_X1 _341_ (
  .A1(_039_),
  .A2(dout[3]),
  .ZN(_077_)
);

NOR2_X2 _342_ (
  .A1(_076_),
  .A2(_077_),
  .ZN(_003_)
);

BUF_X1 _343_ (
  .A(_034_),
  .Z(_078_)
);

NAND2_X1 _344_ (
  .A1(_078_),
  .A2(dout[4]),
  .ZN(_079_)
);

NAND2_X4 _345_ (
  .A1(_062_),
  .A2(_074_),
  .ZN(_080_)
);

INV_X4 _346_ (
  .A(_080_),
  .ZN(_081_)
);

OAI21_X2 _347_ (
  .A(_081_),
  .B1(_055_),
  .B2(_058_),
  .ZN(_082_)
);

NAND2_X2 _348_ (
  .A1(_074_),
  .A2(_275_),
  .ZN(_083_)
);

INV_X1 _349_ (
  .A(_277_),
  .ZN(_084_)
);

NAND2_X2 _350_ (
  .A1(_083_),
  .A2(_084_),
  .ZN(_085_)
);

INV_X1 _351_ (
  .A(_085_),
  .ZN(_086_)
);

NAND2_X2 _352_ (
  .A1(_082_),
  .A2(_086_),
  .ZN(_087_)
);

BUF_X4 _353_ (
  .A(_280_),
  .Z(_088_)
);

XNOR2_X1 _354_ (
  .A(_087_),
  .B(_088_),
  .ZN(_089_)
);

AND2_X2 _355_ (
  .A1(_089_),
  .A2(_037_),
  .ZN(_090_)
);

OAI21_X1 _356_ (
  .A(_039_),
  .B1(_041_),
  .B2(\iq[5] ),
  .ZN(_091_)
);

OAI21_X2 _357_ (
  .A(_079_),
  .B1(_090_),
  .B2(_091_),
  .ZN(_004_)
);

NAND2_X1 _358_ (
  .A1(_078_),
  .A2(dout[5]),
  .ZN(_092_)
);

NAND2_X4 _359_ (
  .A1(_074_),
  .A2(_088_),
  .ZN(_093_)
);

NOR2_X4 _360_ (
  .A1(_072_),
  .A2(_093_),
  .ZN(_094_)
);

NAND2_X2 _361_ (
  .A1(_094_),
  .A2(_045_),
  .ZN(_095_)
);

NAND2_X2 _362_ (
  .A1(_088_),
  .A2(_277_),
  .ZN(_096_)
);

INV_X1 _363_ (
  .A(_279_),
  .ZN(_097_)
);

NAND2_X1 _364_ (
  .A1(_096_),
  .A2(_097_),
  .ZN(_098_)
);

INV_X2 _365_ (
  .A(_098_),
  .ZN(_099_)
);

INV_X2 _366_ (
  .A(_093_),
  .ZN(_100_)
);

NAND2_X2 _367_ (
  .A1(_070_),
  .A2(_100_),
  .ZN(_101_)
);

NAND3_X2 _368_ (
  .A1(_095_),
  .A2(_099_),
  .A3(_101_),
  .ZN(_102_)
);

BUF_X4 _369_ (
  .A(_282_),
  .Z(_103_)
);

XOR2_X2 _370_ (
  .A(_102_),
  .B(_103_),
  .Z(_104_)
);

NOR2_X2 _371_ (
  .A1(_104_),
  .A2(_049_),
  .ZN(_105_)
);

OAI21_X1 _372_ (
  .A(_039_),
  .B1(_041_),
  .B2(\iq[6] ),
  .ZN(_106_)
);

OAI21_X2 _373_ (
  .A(_092_),
  .B1(_105_),
  .B2(_106_),
  .ZN(_005_)
);

NAND2_X4 _374_ (
  .A1(_088_),
  .A2(_103_),
  .ZN(_107_)
);

INV_X4 _375_ (
  .A(_107_),
  .ZN(_108_)
);

NAND3_X2 _376_ (
  .A1(_060_),
  .A2(_081_),
  .A3(_108_),
  .ZN(_109_)
);

NAND2_X1 _377_ (
  .A1(_085_),
  .A2(_108_),
  .ZN(_110_)
);

NAND2_X1 _378_ (
  .A1(_103_),
  .A2(_279_),
  .ZN(_111_)
);

INV_X1 _379_ (
  .A(_281_),
  .ZN(_112_)
);

NAND2_X1 _380_ (
  .A1(_111_),
  .A2(_112_),
  .ZN(_113_)
);

INV_X2 _381_ (
  .A(_113_),
  .ZN(_114_)
);

NAND2_X2 _382_ (
  .A1(_110_),
  .A2(_114_),
  .ZN(_115_)
);

INV_X1 _383_ (
  .A(_115_),
  .ZN(_116_)
);

NAND2_X1 _384_ (
  .A1(_109_),
  .A2(_116_),
  .ZN(_117_)
);

BUF_X4 _385_ (
  .A(_284_),
  .Z(_118_)
);

INV_X1 _386_ (
  .A(_118_),
  .ZN(_119_)
);

NAND2_X1 _387_ (
  .A1(_117_),
  .A2(_119_),
  .ZN(_120_)
);

NAND3_X1 _388_ (
  .A1(_109_),
  .A2(_116_),
  .A3(_118_),
  .ZN(_121_)
);

NAND3_X1 _389_ (
  .A1(_120_),
  .A2(_121_),
  .A3(_041_),
  .ZN(_122_)
);

INV_X1 _390_ (
  .A(\iq[7] ),
  .ZN(_123_)
);

AOI21_X1 _391_ (
  .A(_035_),
  .B1(_049_),
  .B2(_123_),
  .ZN(_124_)
);

NAND2_X1 _392_ (
  .A1(_122_),
  .A2(_124_),
  .ZN(_125_)
);

NAND2_X1 _393_ (
  .A1(_078_),
  .A2(dout[6]),
  .ZN(_126_)
);

NAND2_X1 _394_ (
  .A1(_125_),
  .A2(_126_),
  .ZN(_006_)
);

NAND2_X2 _395_ (
  .A1(_103_),
  .A2(_118_),
  .ZN(_127_)
);

NOR2_X1 _396_ (
  .A1(_093_),
  .A2(_127_),
  .ZN(_128_)
);

NAND2_X2 _397_ (
  .A1(_073_),
  .A2(_128_),
  .ZN(_129_)
);

NAND2_X1 _398_ (
  .A1(_118_),
  .A2(_281_),
  .ZN(_130_)
);

INV_X1 _399_ (
  .A(_283_),
  .ZN(_131_)
);

NAND2_X1 _400_ (
  .A1(_130_),
  .A2(_131_),
  .ZN(_132_)
);

INV_X1 _401_ (
  .A(_132_),
  .ZN(_133_)
);

OAI21_X1 _402_ (
  .A(_133_),
  .B1(_099_),
  .B2(_127_),
  .ZN(_134_)
);

INV_X1 _403_ (
  .A(_134_),
  .ZN(_135_)
);

NAND2_X2 _404_ (
  .A1(_129_),
  .A2(_135_),
  .ZN(_136_)
);

BUF_X4 _405_ (
  .A(_286_),
  .Z(_137_)
);

INV_X1 _406_ (
  .A(_137_),
  .ZN(_138_)
);

NAND2_X1 _407_ (
  .A1(_136_),
  .A2(_138_),
  .ZN(_139_)
);

NAND3_X1 _408_ (
  .A1(_129_),
  .A2(_137_),
  .A3(_135_),
  .ZN(_140_)
);

NAND3_X1 _409_ (
  .A1(_139_),
  .A2(_140_),
  .A3(_041_),
  .ZN(_141_)
);

INV_X1 _410_ (
  .A(\iq[8] ),
  .ZN(_142_)
);

AOI21_X1 _411_ (
  .A(_035_),
  .B1(_049_),
  .B2(_142_),
  .ZN(_143_)
);

NAND2_X1 _412_ (
  .A1(_141_),
  .A2(_143_),
  .ZN(_144_)
);

NAND2_X1 _413_ (
  .A1(_078_),
  .A2(dout[7]),
  .ZN(_145_)
);

NAND2_X1 _414_ (
  .A1(_144_),
  .A2(_145_),
  .ZN(_007_)
);

NAND2_X4 _415_ (
  .A1(_118_),
  .A2(_137_),
  .ZN(_146_)
);

NOR2_X1 _416_ (
  .A1(_107_),
  .A2(_146_),
  .ZN(_147_)
);

NAND2_X2 _417_ (
  .A1(_087_),
  .A2(_147_),
  .ZN(_148_)
);

NAND2_X1 _418_ (
  .A1(_137_),
  .A2(_283_),
  .ZN(_149_)
);

INV_X1 _419_ (
  .A(_285_),
  .ZN(_150_)
);

NAND2_X1 _420_ (
  .A1(_149_),
  .A2(_150_),
  .ZN(_151_)
);

INV_X1 _421_ (
  .A(_151_),
  .ZN(_152_)
);

OAI21_X1 _422_ (
  .A(_152_),
  .B1(_114_),
  .B2(_146_),
  .ZN(_153_)
);

INV_X1 _423_ (
  .A(_153_),
  .ZN(_154_)
);

NAND2_X1 _424_ (
  .A1(_148_),
  .A2(_154_),
  .ZN(_155_)
);

BUF_X4 _425_ (
  .A(_288_),
  .Z(_156_)
);

INV_X1 _426_ (
  .A(_156_),
  .ZN(_157_)
);

NAND2_X1 _427_ (
  .A1(_155_),
  .A2(_157_),
  .ZN(_158_)
);

NAND3_X1 _428_ (
  .A1(_148_),
  .A2(_156_),
  .A3(_154_),
  .ZN(_159_)
);

NAND3_X1 _429_ (
  .A1(_158_),
  .A2(_159_),
  .A3(_041_),
  .ZN(_160_)
);

INV_X1 _430_ (
  .A(\iq[9] ),
  .ZN(_161_)
);

AOI21_X1 _431_ (
  .A(_035_),
  .B1(_049_),
  .B2(_161_),
  .ZN(_162_)
);

NAND2_X1 _432_ (
  .A1(_160_),
  .A2(_162_),
  .ZN(_163_)
);

NAND2_X1 _433_ (
  .A1(_078_),
  .A2(dout[8]),
  .ZN(_164_)
);

NAND2_X1 _434_ (
  .A1(_163_),
  .A2(_164_),
  .ZN(_008_)
);

NAND2_X1 _435_ (
  .A1(_101_),
  .A2(_099_),
  .ZN(_165_)
);

NAND2_X2 _436_ (
  .A1(_137_),
  .A2(_156_),
  .ZN(_166_)
);

NOR2_X2 _437_ (
  .A1(_127_),
  .A2(_166_),
  .ZN(_167_)
);

NAND2_X1 _438_ (
  .A1(_165_),
  .A2(_167_),
  .ZN(_168_)
);

INV_X1 _439_ (
  .A(_166_),
  .ZN(_169_)
);

NAND2_X1 _440_ (
  .A1(_132_),
  .A2(_169_),
  .ZN(_170_)
);

NAND2_X1 _441_ (
  .A1(_156_),
  .A2(_285_),
  .ZN(_171_)
);

INV_X1 _442_ (
  .A(_287_),
  .ZN(_172_)
);

NAND2_X1 _443_ (
  .A1(_171_),
  .A2(_172_),
  .ZN(_173_)
);

INV_X1 _444_ (
  .A(_173_),
  .ZN(_174_)
);

NAND2_X1 _445_ (
  .A1(_170_),
  .A2(_174_),
  .ZN(_175_)
);

INV_X1 _446_ (
  .A(_175_),
  .ZN(_176_)
);

NAND3_X1 _447_ (
  .A1(_094_),
  .A2(_167_),
  .A3(_045_),
  .ZN(_177_)
);

NAND3_X1 _448_ (
  .A1(_168_),
  .A2(_176_),
  .A3(_177_),
  .ZN(_178_)
);

INV_X1 _449_ (
  .A(_290_),
  .ZN(_179_)
);

NAND2_X1 _450_ (
  .A1(_178_),
  .A2(_179_),
  .ZN(_180_)
);

NAND4_X1 _451_ (
  .A1(_168_),
  .A2(_177_),
  .A3(_176_),
  .A4(_290_),
  .ZN(_181_)
);

NAND3_X1 _452_ (
  .A1(_180_),
  .A2(_181_),
  .A3(_041_),
  .ZN(_182_)
);

INV_X1 _453_ (
  .A(\iq[10] ),
  .ZN(_183_)
);

AOI21_X1 _454_ (
  .A(_035_),
  .B1(_049_),
  .B2(_183_),
  .ZN(_184_)
);

NAND2_X1 _455_ (
  .A1(_182_),
  .A2(_184_),
  .ZN(_185_)
);

NAND2_X1 _456_ (
  .A1(_078_),
  .A2(dout[9]),
  .ZN(_186_)
);

NAND2_X1 _457_ (
  .A1(_185_),
  .A2(_186_),
  .ZN(_009_)
);

INV_X2 _458_ (
  .A(_146_),
  .ZN(_187_)
);

NAND2_X4 _459_ (
  .A1(_156_),
  .A2(_290_),
  .ZN(_188_)
);

INV_X2 _460_ (
  .A(_188_),
  .ZN(_189_)
);

NAND2_X2 _461_ (
  .A1(_187_),
  .A2(_189_),
  .ZN(_190_)
);

INV_X1 _462_ (
  .A(_190_),
  .ZN(_191_)
);

NAND2_X2 _463_ (
  .A1(_115_),
  .A2(_191_),
  .ZN(_192_)
);

NAND2_X4 _464_ (
  .A1(_081_),
  .A2(_108_),
  .ZN(_193_)
);

NOR2_X2 _465_ (
  .A1(_193_),
  .A2(_190_),
  .ZN(_194_)
);

NAND2_X2 _466_ (
  .A1(_194_),
  .A2(_060_),
  .ZN(_195_)
);

INV_X1 _467_ (
  .A(_289_),
  .ZN(_196_)
);

OAI21_X1 _468_ (
  .A(_196_),
  .B1(_179_),
  .B2(_172_),
  .ZN(_197_)
);

INV_X1 _469_ (
  .A(_197_),
  .ZN(_198_)
);

NAND2_X1 _470_ (
  .A1(_151_),
  .A2(_189_),
  .ZN(_199_)
);

NAND2_X1 _471_ (
  .A1(_198_),
  .A2(_199_),
  .ZN(_200_)
);

INV_X2 _472_ (
  .A(_200_),
  .ZN(_201_)
);

XNOR2_X1 _473_ (
  .A(\iq[12] ),
  .B(\iq[11] ),
  .ZN(_202_)
);

INV_X1 _474_ (
  .A(_202_),
  .ZN(_203_)
);

NAND4_X1 _475_ (
  .A1(_192_),
  .A2(_195_),
  .A3(_201_),
  .A4(_203_),
  .ZN(_204_)
);

NAND3_X2 _476_ (
  .A1(_192_),
  .A2(_195_),
  .A3(_201_),
  .ZN(_205_)
);

NAND2_X1 _477_ (
  .A1(_205_),
  .A2(_202_),
  .ZN(_206_)
);

NAND3_X1 _478_ (
  .A1(_204_),
  .A2(_206_),
  .A3(_037_),
  .ZN(_207_)
);

INV_X1 _479_ (
  .A(\iq[11] ),
  .ZN(_208_)
);

AOI21_X1 _480_ (
  .A(_035_),
  .B1(_049_),
  .B2(_208_),
  .ZN(_209_)
);

NAND2_X1 _481_ (
  .A1(_207_),
  .A2(_209_),
  .ZN(_210_)
);

NAND2_X1 _482_ (
  .A1(_078_),
  .A2(dout[10]),
  .ZN(_211_)
);

NAND2_X2 _483_ (
  .A1(_210_),
  .A2(_211_),
  .ZN(_010_)
);

BUF_X1 _484_ (
  .A(dstrb),
  .Z(_212_)
);

NOR2_X1 _485_ (
  .A1(_035_),
  .A2(_212_),
  .ZN(_213_)
);

INV_X1 _486_ (
  .A(\dep[0] ),
  .ZN(_214_)
);

AOI21_X1 _487_ (
  .A(_213_),
  .B1(_214_),
  .B2(_078_),
  .ZN(_011_)
);

NAND2_X1 _488_ (
  .A1(_078_),
  .A2(\dep[1] ),
  .ZN(_215_)
);

OAI21_X1 _489_ (
  .A(_215_),
  .B1(_078_),
  .B2(_214_),
  .ZN(_012_)
);

MUX2_X1 _490_ (
  .A(\dep[2] ),
  .B(\dep[1] ),
  .S(_039_),
  .Z(_013_)
);

BUF_X2 _491_ (
  .A(_033_),
  .Z(_216_)
);

MUX2_X1 _492_ (
  .A(\dep[3] ),
  .B(\dep[2] ),
  .S(_216_),
  .Z(_014_)
);

MUX2_X1 _493_ (
  .A(\dep[4] ),
  .B(\dep[3] ),
  .S(_216_),
  .Z(_015_)
);

MUX2_X1 _494_ (
  .A(\dep[5] ),
  .B(\dep[4] ),
  .S(_216_),
  .Z(_016_)
);

MUX2_X1 _495_ (
  .A(\dep[6] ),
  .B(\dep[5] ),
  .S(_033_),
  .Z(_017_)
);

MUX2_X1 _496_ (
  .A(\dep[7] ),
  .B(\dep[6] ),
  .S(_216_),
  .Z(_018_)
);

MUX2_X1 _497_ (
  .A(\dep[8] ),
  .B(\dep[7] ),
  .S(_216_),
  .Z(_019_)
);

MUX2_X1 _498_ (
  .A(\dep[9] ),
  .B(\dep[8] ),
  .S(_216_),
  .Z(_020_)
);

MUX2_X1 _499_ (
  .A(\dep[10] ),
  .B(\dep[9] ),
  .S(_216_),
  .Z(_021_)
);

MUX2_X1 _500_ (
  .A(\dep[11] ),
  .B(\dep[10] ),
  .S(_216_),
  .Z(_022_)
);

MUX2_X1 _501_ (
  .A(\dep[12] ),
  .B(\dep[11] ),
  .S(_216_),
  .Z(_023_)
);

MUX2_X1 _502_ (
  .A(\dep[13] ),
  .B(\dep[12] ),
  .S(_039_),
  .Z(_024_)
);

MUX2_X1 _503_ (
  .A(\dep[14] ),
  .B(\dep[13] ),
  .S(_216_),
  .Z(_025_)
);

MUX2_X1 _504_ (
  .A(douten),
  .B(\dep[14] ),
  .S(_039_),
  .Z(_026_)
);

NAND2_X1 _505_ (
  .A1(_033_),
  .A2(qnt_cnt[0]),
  .ZN(_217_)
);

INV_X1 _506_ (
  .A(_217_),
  .ZN(_218_)
);

NOR2_X1 _507_ (
  .A1(_039_),
  .A2(qnt_cnt[0]),
  .ZN(_219_)
);

NOR3_X1 _508_ (
  .A1(_218_),
  .A2(_219_),
  .A3(_212_),
  .ZN(_027_)
);

NAND2_X1 _509_ (
  .A1(_213_),
  .A2(_292_),
  .ZN(_220_)
);

NAND2_X1 _510_ (
  .A1(_035_),
  .A2(qnt_cnt[1]),
  .ZN(_221_)
);

OAI21_X1 _511_ (
  .A(_220_),
  .B1(_212_),
  .B2(_221_),
  .ZN(_028_)
);

INV_X1 _512_ (
  .A(_291_),
  .ZN(_222_)
);

INV_X1 _513_ (
  .A(qnt_cnt[2]),
  .ZN(_223_)
);

NOR3_X1 _514_ (
  .A1(_034_),
  .A2(_222_),
  .A3(_223_),
  .ZN(_224_)
);

OAI21_X1 _515_ (
  .A(_223_),
  .B1(_034_),
  .B2(_222_),
  .ZN(_225_)
);

INV_X1 _516_ (
  .A(_225_),
  .ZN(_226_)
);

NOR3_X1 _517_ (
  .A1(_224_),
  .A2(_226_),
  .A3(_212_),
  .ZN(_029_)
);

AND3_X2 _518_ (
  .A1(_218_),
  .A2(qnt_cnt[2]),
  .A3(qnt_cnt[1]),
  .ZN(_227_)
);

NAND2_X2 _519_ (
  .A1(_227_),
  .A2(qnt_cnt[3]),
  .ZN(_228_)
);

INV_X1 _520_ (
  .A(_228_),
  .ZN(_229_)
);

NOR2_X1 _521_ (
  .A1(_227_),
  .A2(qnt_cnt[3]),
  .ZN(_230_)
);

NOR3_X1 _522_ (
  .A1(_229_),
  .A2(_230_),
  .A3(_212_),
  .ZN(_030_)
);

AND3_X1 _523_ (
  .A1(_224_),
  .A2(qnt_cnt[3]),
  .A3(qnt_cnt[4]),
  .ZN(_231_)
);

AOI21_X1 _524_ (
  .A(qnt_cnt[4]),
  .B1(_224_),
  .B2(qnt_cnt[3]),
  .ZN(_232_)
);

NOR3_X2 _525_ (
  .A1(_231_),
  .A2(_232_),
  .A3(_212_),
  .ZN(_031_)
);

INV_X1 _526_ (
  .A(qnt_cnt[5]),
  .ZN(_233_)
);

INV_X1 _527_ (
  .A(qnt_cnt[4]),
  .ZN(_234_)
);

OAI21_X1 _528_ (
  .A(_233_),
  .B1(_228_),
  .B2(_234_),
  .ZN(_235_)
);

INV_X1 _529_ (
  .A(_235_),
  .ZN(_236_)
);

NOR3_X1 _530_ (
  .A1(_228_),
  .A2(_234_),
  .A3(_233_),
  .ZN(_237_)
);

NOR3_X2 _531_ (
  .A1(_236_),
  .A2(_237_),
  .A3(_212_),
  .ZN(_032_)
);

HA_X1 _532_ (
  .A(\iq[1] ),
  .B(\iq[12] ),
  .CO(_271_),
  .S(_272_)
);

HA_X1 _533_ (
  .A(\iq[2] ),
  .B(\iq[12] ),
  .CO(_273_),
  .S(_274_)
);

HA_X1 _534_ (
  .A(\iq[3] ),
  .B(\iq[12] ),
  .CO(_275_),
  .S(_276_)
);

HA_X1 _535_ (
  .A(\iq[4] ),
  .B(\iq[12] ),
  .CO(_277_),
  .S(_278_)
);

HA_X1 _536_ (
  .A(\iq[5] ),
  .B(\iq[12] ),
  .CO(_279_),
  .S(_280_)
);

HA_X1 _537_ (
  .A(\iq[6] ),
  .B(\iq[12] ),
  .CO(_281_),
  .S(_282_)
);

HA_X1 _538_ (
  .A(\iq[7] ),
  .B(\iq[12] ),
  .CO(_283_),
  .S(_284_)
);

HA_X1 _539_ (
  .A(\iq[8] ),
  .B(\iq[12] ),
  .CO(_285_),
  .S(_286_)
);

HA_X1 _540_ (
  .A(\iq[9] ),
  .B(\iq[12] ),
  .CO(_287_),
  .S(_288_)
);

HA_X1 _541_ (
  .A(\iq[10] ),
  .B(\iq[12] ),
  .CO(_289_),
  .S(_290_)
);

HA_X1 _542_ (
  .A(qnt_cnt[0]),
  .B(qnt_cnt[1]),
  .CO(_291_),
  .S(_292_)
);

LOGIC0_X1 _543_ (
  .Z(_293_)
);

DFFR_X1 \dep[0]$_DFFE_PN0P_  (
  .D(_011_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[0] ),
  .QN(_259_)
);

DFFR_X1 \dep[10]$_DFFE_PN0P_  (
  .D(_021_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[10] ),
  .QN(_249_)
);

DFFR_X1 \dep[11]$_DFFE_PN0P_  (
  .D(_022_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[11] ),
  .QN(_248_)
);

DFFR_X1 \dep[12]$_DFFE_PN0P_  (
  .D(_023_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[12] ),
  .QN(_247_)
);

DFFR_X1 \dep[13]$_DFFE_PN0P_  (
  .D(_024_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[13] ),
  .QN(_246_)
);

DFFR_X1 \dep[14]$_DFFE_PN0P_  (
  .D(_025_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[14] ),
  .QN(_245_)
);

DFFR_X1 \dep[1]$_DFFE_PN0P_  (
  .D(_012_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[1] ),
  .QN(_258_)
);

DFFR_X1 \dep[2]$_DFFE_PN0P_  (
  .D(_013_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[2] ),
  .QN(_257_)
);

DFFR_X1 \dep[3]$_DFFE_PN0P_  (
  .D(_014_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[3] ),
  .QN(_256_)
);

DFFR_X1 \dep[4]$_DFFE_PN0P_  (
  .D(_015_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[4] ),
  .QN(_255_)
);

DFFR_X1 \dep[5]$_DFFE_PN0P_  (
  .D(_016_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[5] ),
  .QN(_254_)
);

DFFR_X1 \dep[6]$_DFFE_PN0P_  (
  .D(_017_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[6] ),
  .QN(_253_)
);

DFFR_X1 \dep[7]$_DFFE_PN0P_  (
  .D(_018_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[7] ),
  .QN(_252_)
);

DFFR_X1 \dep[8]$_DFFE_PN0P_  (
  .D(_019_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[8] ),
  .QN(_251_)
);

DFFR_X1 \dep[9]$_DFFE_PN0P_  (
  .D(_020_),
  .RN(rst),
  .CK(clk),
  .Q(\dep[9] ),
  .QN(_250_)
);

\$paramod\div_su\z_width=s32'00000000000000000000000000011000  divider (
  .clk(clk),
  .ena(ena),
  .z({din[11], din[11], din[11], din[11], din[11], din[11], din[11], din[11], din[11], din[11], din[11], din[11], din}),
  .d({_293_, _293_, _293_, _293_, qnt_val}),
  .q({\iq[12] , \iq[11] , \iq[10] , \iq[9] , \iq[8] , \iq[7] , \iq[6] , \iq[5] , \iq[4] , \iq[3] , \iq[2] , \iq[1] , \iq[0] })
);

DFF_X1 \dout[0]$_DFFE_PP_  (
  .D(_000_),
  .CK(clk),
  .Q(dout[0]),
  .QN(_270_)
);

DFF_X1 \dout[10]$_DFFE_PP_  (
  .D(_010_),
  .CK(clk),
  .Q(dout[10]),
  .QN(_260_)
);

DFF_X1 \dout[1]$_DFFE_PP_  (
  .D(_001_),
  .CK(clk),
  .Q(dout[1]),
  .QN(_269_)
);

DFF_X1 \dout[2]$_DFFE_PP_  (
  .D(_002_),
  .CK(clk),
  .Q(dout[2]),
  .QN(_268_)
);

DFF_X1 \dout[3]$_DFFE_PP_  (
  .D(_003_),
  .CK(clk),
  .Q(dout[3]),
  .QN(_267_)
);

DFF_X1 \dout[4]$_DFFE_PP_  (
  .D(_004_),
  .CK(clk),
  .Q(dout[4]),
  .QN(_266_)
);

DFF_X1 \dout[5]$_DFFE_PP_  (
  .D(_005_),
  .CK(clk),
  .Q(dout[5]),
  .QN(_265_)
);

DFF_X1 \dout[6]$_DFFE_PP_  (
  .D(_006_),
  .CK(clk),
  .Q(dout[6]),
  .QN(_264_)
);

DFF_X1 \dout[7]$_DFFE_PP_  (
  .D(_007_),
  .CK(clk),
  .Q(dout[7]),
  .QN(_263_)
);

DFF_X1 \dout[8]$_DFFE_PP_  (
  .D(_008_),
  .CK(clk),
  .Q(dout[8]),
  .QN(_262_)
);

DFF_X1 \dout[9]$_DFFE_PP_  (
  .D(_009_),
  .CK(clk),
  .Q(dout[9]),
  .QN(_261_)
);

DFFR_X1 douten$_DFFE_PN0P_ (
  .D(_026_),
  .RN(rst),
  .CK(clk),
  .Q(douten),
  .QN(_244_)
);

DFFR_X1 \qnt_cnt[0]$_DFFE_PN0P_  (
  .D(_027_),
  .RN(rst),
  .CK(clk),
  .Q(qnt_cnt[0]),
  .QN(_243_)
);

DFFR_X1 \qnt_cnt[1]$_DFFE_PN0P_  (
  .D(_028_),
  .RN(rst),
  .CK(clk),
  .Q(qnt_cnt[1]),
  .QN(_242_)
);

DFFR_X1 \qnt_cnt[2]$_DFFE_PN0P_  (
  .D(_029_),
  .RN(rst),
  .CK(clk),
  .Q(qnt_cnt[2]),
  .QN(_241_)
);

DFFR_X1 \qnt_cnt[3]$_DFFE_PN0P_  (
  .D(_030_),
  .RN(rst),
  .CK(clk),
  .Q(qnt_cnt[3]),
  .QN(_240_)
);

DFFR_X1 \qnt_cnt[4]$_DFFE_PN0P_  (
  .D(_031_),
  .RN(rst),
  .CK(clk),
  .Q(qnt_cnt[4]),
  .QN(_239_)
);

DFFR_X1 \qnt_cnt[5]$_DFFE_PN0P_  (
  .D(_032_),
  .RN(rst),
  .CK(clk),
  .Q(qnt_cnt[5]),
  .QN(_238_)
);
endmodule //jpeg_qnr

module \$paramod$bae1c4187f9f11528499493f4465458a121f3954\dctub (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout0, output [11:0] dout1,
 output [11:0] dout2, output [11:0] dout3, output [11:0] dout4, output [11:0] dout5, output [11:0] dout6,
 output [11:0] dout7);
\$paramod$2da196d8114b669d4bb3858ca0a91434452576e0\dctu  dct_unit_0 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout0)
);

\$paramod$a5796bae454a3870edf919a9404bde7ca4192701\dctu  dct_unit_1 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout1)
);

\$paramod$eb0441514cb1002bdcaf5201d3067d7bd1bbd3e9\dctu  dct_unit_2 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout2)
);

\$paramod$e9d96eb14c78f030ece167996f154f4849a68288\dctu  dct_unit_3 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout3)
);

\$paramod$2ce29d501700894abc3f54c094daafc2d8c2c211\dctu  dct_unit_4 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout4)
);

\$paramod$11fa2caec0040cf5bdd9aac167c50c8009d1fe68\dctu  dct_unit_5 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout5)
);

\$paramod$bd585d540938973e77d9fdfafe68a3c54bf55cb8\dctu  dct_unit_6 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout6)
);

\$paramod$94a1b10314722615b96d6c8f661cbb82ecebf320\dctu  dct_unit_7 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout7)
);
endmodule //$paramod$bae1c4187f9f11528499493f4465458a121f3954\dctub

module \$paramod$10132426324c91f74f0d67bb39d4db77efb06075\dctub (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout0, output [11:0] dout1,
 output [11:0] dout2, output [11:0] dout3, output [11:0] dout4, output [11:0] dout5, output [11:0] dout6,
 output [11:0] dout7);
\$paramod$53ab2e60687d01e7461fdffe1d34a14bacda6928\dctu  dct_unit_0 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout0)
);

\$paramod$99c498a68fd2923ba65be259bfb6e7d8309d79f4\dctu  dct_unit_1 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout1)
);

\$paramod$f5bb6813249a03e2893277297591ec050ac518dc\dctu  dct_unit_2 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout2)
);

\$paramod$696f85e1ea63d2b5ad7171a625fd3b51a665057d\dctu  dct_unit_3 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout3)
);

\$paramod$8f6708f3156f3d6d195809cddd67c9b8c08cd488\dctu  dct_unit_4 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout4)
);

\$paramod$e2471d3acfddfd8f107137e4952b02d9e7720f44\dctu  dct_unit_5 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout5)
);

\$paramod$9e8342fceac8003655f9e71995b4fdeb8565fbe5\dctu  dct_unit_6 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout6)
);

\$paramod$0f96740a02eb44c944b68d6b495a8cce162f1249\dctu  dct_unit_7 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout7)
);
endmodule //$paramod$10132426324c91f74f0d67bb39d4db77efb06075\dctub

module \$paramod$0b8c49989cad027b3dfd23a8cec031b2f9a47f64\dctub (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout0, output [11:0] dout1,
 output [11:0] dout2, output [11:0] dout3, output [11:0] dout4, output [11:0] dout5, output [11:0] dout6,
 output [11:0] dout7);
\$paramod$3b47752d19f391915a818678f43c9a51f524cc48\dctu  dct_unit_0 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout0)
);

\$paramod$b266e2f77428397c53d4afd55bef1da32efe03d9\dctu  dct_unit_1 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout1)
);

\$paramod$f06914ec453560c29e1738d8a2be788b84af024b\dctu  dct_unit_2 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout2)
);

\$paramod$a184ef4c0e9b8e48eac4b335f6b36fd82c0c32d3\dctu  dct_unit_3 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout3)
);

\$paramod$6be19b0824fdb8c44e931702b04949b1ae101a34\dctu  dct_unit_4 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout4)
);

\$paramod$1b119bd029c81aaa2221a23d15ab3b6b02f6efee\dctu  dct_unit_5 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout5)
);

\$paramod$9fe6c97945bcc341eadabee9cbdea0f75515e5c3\dctu  dct_unit_6 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout6)
);

\$paramod$44a044575968c599376fc32b4d9ee49faea5711d\dctu  dct_unit_7 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout7)
);
endmodule //$paramod$0b8c49989cad027b3dfd23a8cec031b2f9a47f64\dctub

module \$paramod$08d1c923a0daedefe47ae23865eeb002e5733497\dctub (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout0, output [11:0] dout1,
 output [11:0] dout2, output [11:0] dout3, output [11:0] dout4, output [11:0] dout5, output [11:0] dout6,
 output [11:0] dout7);
\$paramod$e6bd937dcb54fb0697fee40c5f9824ba6fd53538\dctu  dct_unit_0 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout0)
);

\$paramod$da3415da01ee30cd3fa431ef7b8104a7c6ed9a24\dctu  dct_unit_1 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout1)
);

\$paramod$b53123087aafc52fe604e5dcf6b6b1b8d73b2231\dctu  dct_unit_2 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout2)
);

\$paramod$4dc5718e86f31fe555f7d39cf5ab7078c09f577a\dctu  dct_unit_3 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout3)
);

\$paramod$fa41e4d02884503da5d6c381e868b8c261424a31\dctu  dct_unit_4 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout4)
);

\$paramod$826cb5d104d530340b1f58495d2410742b2c32fe\dctu  dct_unit_5 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout5)
);

\$paramod$88a8287894fa5d106cca0ce24429339f4a2785a9\dctu  dct_unit_6 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout6)
);

\$paramod$0c5a5bd6be4ed818deaac08b02afbddb6897ffee\dctu  dct_unit_7 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout7)
);
endmodule //$paramod$08d1c923a0daedefe47ae23865eeb002e5733497\dctub

module \$paramod$5da4b737faccfde9a093da147c1f0b2523b6c7dd\dctub (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout0, output [11:0] dout1,
 output [11:0] dout2, output [11:0] dout3, output [11:0] dout4, output [11:0] dout5, output [11:0] dout6,
 output [11:0] dout7);
\$paramod$d348381a5c8d7c369f0c055d305d608d67b77e86\dctu  dct_unit_0 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout0)
);

\$paramod$29130e85acc43116076719ea36da8d59b7490cc4\dctu  dct_unit_1 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout1)
);

\$paramod$32a02d514417e24bb09b7885b9c053483ac7784d\dctu  dct_unit_2 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout2)
);

\$paramod$9beaa443332981731011e314e41ebdfa5267d059\dctu  dct_unit_3 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout3)
);

\$paramod$fa85f450a22557b2687ca86acb15721a7fddf8e7\dctu  dct_unit_4 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout4)
);

\$paramod$5778094f610ca183dd46956f589e4ea513d2316c\dctu  dct_unit_5 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout5)
);

\$paramod$cf6677181b8958913bf11288905dc7e6338a7bf5\dctu  dct_unit_6 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout6)
);

\$paramod$4895890460618319d2e2de05b5a45e21ba9e3f8b\dctu  dct_unit_7 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout7)
);
endmodule //$paramod$5da4b737faccfde9a093da147c1f0b2523b6c7dd\dctub

module \$paramod$47ef26d4334fc5e08bebdeabebd3eea4dff44a0a\dctub (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout0, output [11:0] dout1,
 output [11:0] dout2, output [11:0] dout3, output [11:0] dout4, output [11:0] dout5, output [11:0] dout6,
 output [11:0] dout7);
\$paramod$f1b01728a98736f8d413a71bd9a7600c5a6961e3\dctu  dct_unit_0 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout0)
);

\$paramod$04fdc4f446e06e0744e44efd615d1158fec3aeb8\dctu  dct_unit_1 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout1)
);

\$paramod$a523c923d4f86f07f4e81f5d8b04b352dfcc17be\dctu  dct_unit_2 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout2)
);

\$paramod$c4f8cc56c0ef9356356d2a98d35862f209dd307b\dctu  dct_unit_3 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout3)
);

\$paramod$adcdc49d3fc5249816d353bb65629f56cf0927d3\dctu  dct_unit_4 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout4)
);

\$paramod$bfc28a02cfebf191b4a982c9147f38f65a3f3469\dctu  dct_unit_5 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout5)
);

\$paramod$7911a3968b23dded19efefb86cf26bb44e3a7781\dctu  dct_unit_6 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout6)
);

\$paramod$785fe1ea8cdf428cbeb2f89081ee68c33feb7da2\dctu  dct_unit_7 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout7)
);
endmodule //$paramod$47ef26d4334fc5e08bebdeabebd3eea4dff44a0a\dctub

module \$paramod$302a2dacc76057b68e5fd92243d54f2e7b35812d\dctub (input clk, input ena,
 input ddgo, input [2:0] x, input [2:0] y, input [8:1] ddin, output [11:0] dout0, output [11:0] dout1,
 output [11:0] dout2, output [11:0] dout3, output [11:0] dout4, output [11:0] dout5, output [11:0] dout6,
 output [11:0] dout7);
\$paramod$141303f1e6ff0436e3fa44dd8e1d8f51afed9a78\dctu  dct_unit_0 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout0)
);

\$paramod$16cad72ebc555f93621a2c70f423f14f85bbeb07\dctu  dct_unit_1 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout1)
);

\$paramod$a8d3b7b4edaf7d596a54a187c8ed4a9561fa625a\dctu  dct_unit_2 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout2)
);

\$paramod$56b31b71c3bccc1fb1f134779b3bdd5ab1b461c7\dctu  dct_unit_3 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout3)
);

\$paramod$141b5017b00a41bd6bcdd772ef8ad836aaf4019f\dctu  dct_unit_4 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout4)
);

\$paramod$37cd075c9fa8b3a4872c05f999800e89bc604dc4\dctu  dct_unit_5 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout5)
);

\$paramod$26ce9ce45d1136272d6a188b0b22329681d6199b\dctu  dct_unit_6 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout6)
);

\$paramod$ca051f171e86125a3bcf4bd090f5be774b98c04e\dctu  dct_unit_7 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x(x),
  .y(y),
  .ddin(ddin),
  .dout(dout7)
);
endmodule //$paramod$302a2dacc76057b68e5fd92243d54f2e7b35812d\dctub

module \$paramod$849c8591669cf197b80ef99050b300773b555aae\dct (input clk, input ena,
 input rst, input dstrb, input [8:1] din, output [12:1] dout_00, output [12:1] dout_01,
 output [12:1] dout_02, output [12:1] dout_03, output [12:1] dout_04, output [12:1] dout_05,
 output [12:1] dout_06, output [12:1] dout_07, output [12:1] dout_10, output [12:1] dout_11,
 output [12:1] dout_12, output [12:1] dout_13, output [12:1] dout_14, output [12:1] dout_15,
 output [12:1] dout_16, output [12:1] dout_17, output [12:1] dout_20, output [12:1] dout_21,
 output [12:1] dout_22, output [12:1] dout_23, output [12:1] dout_24, output [12:1] dout_25,
 output [12:1] dout_26, output [12:1] dout_27, output [12:1] dout_30, output [12:1] dout_31,
 output [12:1] dout_32, output [12:1] dout_33, output [12:1] dout_34, output [12:1] dout_35,
 output [12:1] dout_36, output [12:1] dout_37, output [12:1] dout_40, output [12:1] dout_41,
 output [12:1] dout_42, output [12:1] dout_43, output [12:1] dout_44, output [12:1] dout_45,
 output [12:1] dout_46, output [12:1] dout_47, output [12:1] dout_50, output [12:1] dout_51,
 output [12:1] dout_52, output [12:1] dout_53, output [12:1] dout_54, output [12:1] dout_55,
 output [12:1] dout_56, output [12:1] dout_57, output [12:1] dout_60, output [12:1] dout_61,
 output [12:1] dout_62, output [12:1] dout_63, output [12:1] dout_64, output [12:1] dout_65,
 output [12:1] dout_66, output [12:1] dout_67, output [12:1] dout_70, output [12:1] dout_71,
 output [12:1] dout_72, output [12:1] dout_73, output [12:1] dout_74, output [12:1] dout_75,
 output [12:1] dout_76, output [12:1] dout_77, output douten);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire ddcnt;
wire dddcnt;
wire ddgo;
wire \ddin[1] ;
wire \ddin[2] ;
wire \ddin[3] ;
wire \ddin[4] ;
wire \ddin[5] ;
wire \ddin[6] ;
wire \ddin[7] ;
wire \ddin[8] ;
wire dgo;
wire go;
wire \sample_cnt[0] ;
wire \sample_cnt[1] ;
wire \sample_cnt[2] ;
wire \sample_cnt[3] ;
wire \sample_cnt[4] ;
wire \sample_cnt[5] ;

BUF_X4 _085_ (
  .A(ena),
  .Z(_023_)
);

BUF_X4 _086_ (
  .A(\sample_cnt[3] ),
  .Z(_024_)
);

BUF_X4 _087_ (
  .A(\sample_cnt[2] ),
  .Z(_025_)
);

NAND3_X4 _088_ (
  .A1(_024_),
  .A2(_025_),
  .A3(_083_),
  .ZN(_026_)
);

NAND2_X1 _089_ (
  .A1(\sample_cnt[5] ),
  .A2(\sample_cnt[4] ),
  .ZN(_027_)
);

OAI21_X4 _090_ (
  .A(_023_),
  .B1(_026_),
  .B2(_027_),
  .ZN(_028_)
);

BUF_X1 _091_ (
  .A(dstrb),
  .Z(_029_)
);

NAND2_X2 _092_ (
  .A1(_029_),
  .A2(_023_),
  .ZN(_030_)
);

NAND2_X4 _093_ (
  .A1(_028_),
  .A2(_030_),
  .ZN(_031_)
);

INV_X1 _094_ (
  .A(_029_),
  .ZN(_032_)
);

INV_X1 _095_ (
  .A(\sample_cnt[0] ),
  .ZN(_033_)
);

NAND3_X1 _096_ (
  .A1(_031_),
  .A2(_032_),
  .A3(_033_),
  .ZN(_034_)
);

NAND3_X1 _097_ (
  .A1(_028_),
  .A2(\sample_cnt[0] ),
  .A3(_030_),
  .ZN(_035_)
);

NAND2_X1 _098_ (
  .A1(_034_),
  .A2(_035_),
  .ZN(_000_)
);

NAND3_X1 _099_ (
  .A1(_028_),
  .A2(\sample_cnt[1] ),
  .A3(_030_),
  .ZN(_036_)
);

NAND2_X1 _100_ (
  .A1(_032_),
  .A2(_084_),
  .ZN(_037_)
);

OAI21_X1 _101_ (
  .A(_036_),
  .B1(_028_),
  .B2(_037_),
  .ZN(_001_)
);

OR2_X1 _102_ (
  .A1(_083_),
  .A2(_025_),
  .ZN(_038_)
);

NAND2_X1 _103_ (
  .A1(_025_),
  .A2(_083_),
  .ZN(_039_)
);

NAND3_X1 _104_ (
  .A1(_038_),
  .A2(_032_),
  .A3(_039_),
  .ZN(_040_)
);

INV_X1 _105_ (
  .A(_040_),
  .ZN(_041_)
);

NAND2_X1 _106_ (
  .A1(_031_),
  .A2(_041_),
  .ZN(_042_)
);

INV_X1 _107_ (
  .A(_025_),
  .ZN(_043_)
);

OAI21_X2 _108_ (
  .A(_042_),
  .B1(_043_),
  .B2(_031_),
  .ZN(_002_)
);

NAND3_X2 _109_ (
  .A1(_025_),
  .A2(\sample_cnt[0] ),
  .A3(\sample_cnt[1] ),
  .ZN(_044_)
);

XNOR2_X1 _110_ (
  .A(_044_),
  .B(_024_),
  .ZN(_045_)
);

NAND3_X1 _111_ (
  .A1(_031_),
  .A2(_032_),
  .A3(_045_),
  .ZN(_046_)
);

NAND3_X1 _112_ (
  .A1(_028_),
  .A2(_024_),
  .A3(_030_),
  .ZN(_047_)
);

NAND2_X1 _113_ (
  .A1(_046_),
  .A2(_047_),
  .ZN(_003_)
);

NAND2_X1 _114_ (
  .A1(_024_),
  .A2(\sample_cnt[4] ),
  .ZN(_048_)
);

OR2_X1 _115_ (
  .A1(_048_),
  .A2(_039_),
  .ZN(_049_)
);

INV_X1 _116_ (
  .A(\sample_cnt[4] ),
  .ZN(_050_)
);

AOI21_X1 _117_ (
  .A(_029_),
  .B1(_026_),
  .B2(_050_),
  .ZN(_051_)
);

NAND3_X1 _118_ (
  .A1(_031_),
  .A2(_049_),
  .A3(_051_),
  .ZN(_052_)
);

NAND3_X1 _119_ (
  .A1(_028_),
  .A2(\sample_cnt[4] ),
  .A3(_030_),
  .ZN(_053_)
);

NAND2_X1 _120_ (
  .A1(_052_),
  .A2(_053_),
  .ZN(_004_)
);

NOR2_X1 _121_ (
  .A1(_044_),
  .A2(_048_),
  .ZN(_054_)
);

AOI21_X1 _122_ (
  .A(_029_),
  .B1(_054_),
  .B2(\sample_cnt[5] ),
  .ZN(_055_)
);

OR2_X1 _123_ (
  .A1(_054_),
  .A2(\sample_cnt[5] ),
  .ZN(_056_)
);

NAND3_X1 _124_ (
  .A1(_055_),
  .A2(_031_),
  .A3(_056_),
  .ZN(_057_)
);

NAND3_X1 _125_ (
  .A1(_028_),
  .A2(\sample_cnt[5] ),
  .A3(_030_),
  .ZN(_058_)
);

NAND2_X1 _126_ (
  .A1(_057_),
  .A2(_058_),
  .ZN(_005_)
);

BUF_X4 _127_ (
  .A(_023_),
  .Z(_059_)
);

NAND2_X1 _128_ (
  .A1(_059_),
  .A2(ddcnt),
  .ZN(_060_)
);

INV_X1 _129_ (
  .A(douten),
  .ZN(_061_)
);

OAI22_X1 _130_ (
  .A1(_060_),
  .A2(dddcnt),
  .B1(_061_),
  .B2(_059_),
  .ZN(_006_)
);

INV_X1 _131_ (
  .A(go),
  .ZN(_062_)
);

OAI21_X1 _132_ (
  .A(_030_),
  .B1(_059_),
  .B2(_062_),
  .ZN(_007_)
);

NOR2_X1 _133_ (
  .A1(_059_),
  .A2(dgo),
  .ZN(_020_)
);

AOI21_X1 _134_ (
  .A(_020_),
  .B1(_062_),
  .B2(_059_),
  .ZN(_008_)
);

MUX2_X1 _135_ (
  .A(ddgo),
  .B(dgo),
  .S(_023_),
  .Z(_009_)
);

OR2_X1 _136_ (
  .A1(ddcnt),
  .A2(_023_),
  .ZN(_021_)
);

AND2_X1 _137_ (
  .A1(_028_),
  .A2(_021_),
  .ZN(_010_)
);

INV_X1 _138_ (
  .A(dddcnt),
  .ZN(_022_)
);

OAI21_X1 _139_ (
  .A(_060_),
  .B1(_059_),
  .B2(_022_),
  .ZN(_011_)
);

MUX2_X1 _140_ (
  .A(\ddin[1] ),
  .B(din[1]),
  .S(_023_),
  .Z(_012_)
);

MUX2_X1 _141_ (
  .A(\ddin[2] ),
  .B(din[2]),
  .S(_059_),
  .Z(_013_)
);

MUX2_X1 _142_ (
  .A(\ddin[3] ),
  .B(din[3]),
  .S(_059_),
  .Z(_014_)
);

MUX2_X1 _143_ (
  .A(\ddin[4] ),
  .B(din[4]),
  .S(_059_),
  .Z(_015_)
);

MUX2_X1 _144_ (
  .A(\ddin[5] ),
  .B(din[5]),
  .S(_023_),
  .Z(_016_)
);

MUX2_X1 _145_ (
  .A(\ddin[6] ),
  .B(din[6]),
  .S(_023_),
  .Z(_017_)
);

MUX2_X1 _146_ (
  .A(\ddin[7] ),
  .B(din[7]),
  .S(_059_),
  .Z(_018_)
);

MUX2_X1 _147_ (
  .A(\ddin[8] ),
  .B(din[8]),
  .S(_023_),
  .Z(_019_)
);

HA_X1 _148_ (
  .A(\sample_cnt[0] ),
  .B(\sample_cnt[1] ),
  .CO(_083_),
  .S(_084_)
);

\$paramod$f79433e3440244ebaeb06fcd795abd5555024789\dctub  dct_block_0 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x({\sample_cnt[2] , \sample_cnt[1] , \sample_cnt[0] }),
  .y({\sample_cnt[5] , \sample_cnt[4] , \sample_cnt[3] }),
  .ddin({\ddin[8] , \ddin[7] , \ddin[6] , \ddin[5] , \ddin[4] , \ddin[3] , \ddin[2] , \ddin[1] }),
  .dout0(dout_00),
  .dout1(dout_01),
  .dout2(dout_02),
  .dout3(dout_03),
  .dout4(dout_04),
  .dout5(dout_05),
  .dout6(dout_06),
  .dout7(dout_07)
);

\$paramod$10132426324c91f74f0d67bb39d4db77efb06075\dctub  dct_block_1 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x({\sample_cnt[2] , \sample_cnt[1] , \sample_cnt[0] }),
  .y({\sample_cnt[5] , \sample_cnt[4] , \sample_cnt[3] }),
  .ddin({\ddin[8] , \ddin[7] , \ddin[6] , \ddin[5] , \ddin[4] , \ddin[3] , \ddin[2] , \ddin[1] }),
  .dout0(dout_10),
  .dout1(dout_11),
  .dout2(dout_12),
  .dout3(dout_13),
  .dout4(dout_14),
  .dout5(dout_15),
  .dout6(dout_16),
  .dout7(dout_17)
);

\$paramod$08d1c923a0daedefe47ae23865eeb002e5733497\dctub  dct_block_2 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x({\sample_cnt[2] , \sample_cnt[1] , \sample_cnt[0] }),
  .y({\sample_cnt[5] , \sample_cnt[4] , \sample_cnt[3] }),
  .ddin({\ddin[8] , \ddin[7] , \ddin[6] , \ddin[5] , \ddin[4] , \ddin[3] , \ddin[2] , \ddin[1] }),
  .dout0(dout_20),
  .dout1(dout_21),
  .dout2(dout_22),
  .dout3(dout_23),
  .dout4(dout_24),
  .dout5(dout_25),
  .dout6(dout_26),
  .dout7(dout_27)
);

\$paramod$302a2dacc76057b68e5fd92243d54f2e7b35812d\dctub  dct_block_3 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x({\sample_cnt[2] , \sample_cnt[1] , \sample_cnt[0] }),
  .y({\sample_cnt[5] , \sample_cnt[4] , \sample_cnt[3] }),
  .ddin({\ddin[8] , \ddin[7] , \ddin[6] , \ddin[5] , \ddin[4] , \ddin[3] , \ddin[2] , \ddin[1] }),
  .dout0(dout_30),
  .dout1(dout_31),
  .dout2(dout_32),
  .dout3(dout_33),
  .dout4(dout_34),
  .dout5(dout_35),
  .dout6(dout_36),
  .dout7(dout_37)
);

\$paramod$0b8c49989cad027b3dfd23a8cec031b2f9a47f64\dctub  dct_block_4 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x({\sample_cnt[2] , \sample_cnt[1] , \sample_cnt[0] }),
  .y({\sample_cnt[5] , \sample_cnt[4] , \sample_cnt[3] }),
  .ddin({\ddin[8] , \ddin[7] , \ddin[6] , \ddin[5] , \ddin[4] , \ddin[3] , \ddin[2] , \ddin[1] }),
  .dout0(dout_40),
  .dout1(dout_41),
  .dout2(dout_42),
  .dout3(dout_43),
  .dout4(dout_44),
  .dout5(dout_45),
  .dout6(dout_46),
  .dout7(dout_47)
);

\$paramod$47ef26d4334fc5e08bebdeabebd3eea4dff44a0a\dctub  dct_block_5 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x({\sample_cnt[2] , \sample_cnt[1] , \sample_cnt[0] }),
  .y({\sample_cnt[5] , \sample_cnt[4] , \sample_cnt[3] }),
  .ddin({\ddin[8] , \ddin[7] , \ddin[6] , \ddin[5] , \ddin[4] , \ddin[3] , \ddin[2] , \ddin[1] }),
  .dout0(dout_50),
  .dout1(dout_51),
  .dout2(dout_52),
  .dout3(dout_53),
  .dout4(dout_54),
  .dout5(dout_55),
  .dout6(dout_56),
  .dout7(dout_57)
);

\$paramod$bae1c4187f9f11528499493f4465458a121f3954\dctub  dct_block_6 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x({\sample_cnt[2] , \sample_cnt[1] , \sample_cnt[0] }),
  .y({\sample_cnt[5] , \sample_cnt[4] , \sample_cnt[3] }),
  .ddin({\ddin[8] , \ddin[7] , \ddin[6] , \ddin[5] , \ddin[4] , \ddin[3] , \ddin[2] , \ddin[1] }),
  .dout0(dout_60),
  .dout1(dout_61),
  .dout2(dout_62),
  .dout3(dout_63),
  .dout4(dout_64),
  .dout5(dout_65),
  .dout6(dout_66),
  .dout7(dout_67)
);

\$paramod$5da4b737faccfde9a093da147c1f0b2523b6c7dd\dctub  dct_block_7 (
  .clk(clk),
  .ena(ena),
  .ddgo(ddgo),
  .x({\sample_cnt[2] , \sample_cnt[1] , \sample_cnt[0] }),
  .y({\sample_cnt[5] , \sample_cnt[4] , \sample_cnt[3] }),
  .ddin({\ddin[8] , \ddin[7] , \ddin[6] , \ddin[5] , \ddin[4] , \ddin[3] , \ddin[2] , \ddin[1] }),
  .dout0(dout_70),
  .dout1(dout_71),
  .dout2(dout_72),
  .dout3(dout_73),
  .dout4(dout_74),
  .dout5(dout_75),
  .dout6(dout_76),
  .dout7(dout_77)
);

DFFS_X1 ddcnt$_DFFE_PN1P_ (
  .D(_010_),
  .SN(rst),
  .CK(clk),
  .Q(ddcnt),
  .QN(_072_)
);

DFFS_X1 dddcnt$_DFFE_PN1P_ (
  .D(_011_),
  .SN(rst),
  .CK(clk),
  .Q(dddcnt),
  .QN(_071_)
);

DFFR_X1 ddgo$_DFFE_PN0P_ (
  .D(_009_),
  .RN(rst),
  .CK(clk),
  .Q(ddgo),
  .QN(_073_)
);

DFFR_X1 \ddin[0]$_DFFE_PN0P_  (
  .D(_012_),
  .RN(rst),
  .CK(clk),
  .Q(\ddin[1] ),
  .QN(_070_)
);

DFFR_X1 \ddin[1]$_DFFE_PN0P_  (
  .D(_013_),
  .RN(rst),
  .CK(clk),
  .Q(\ddin[2] ),
  .QN(_069_)
);

DFFR_X1 \ddin[2]$_DFFE_PN0P_  (
  .D(_014_),
  .RN(rst),
  .CK(clk),
  .Q(\ddin[3] ),
  .QN(_068_)
);

DFFR_X1 \ddin[3]$_DFFE_PN0P_  (
  .D(_015_),
  .RN(rst),
  .CK(clk),
  .Q(\ddin[4] ),
  .QN(_067_)
);

DFFR_X1 \ddin[4]$_DFFE_PN0P_  (
  .D(_016_),
  .RN(rst),
  .CK(clk),
  .Q(\ddin[5] ),
  .QN(_066_)
);

DFFR_X1 \ddin[5]$_DFFE_PN0P_  (
  .D(_017_),
  .RN(rst),
  .CK(clk),
  .Q(\ddin[6] ),
  .QN(_065_)
);

DFFR_X1 \ddin[6]$_DFFE_PN0P_  (
  .D(_018_),
  .RN(rst),
  .CK(clk),
  .Q(\ddin[7] ),
  .QN(_064_)
);

DFFR_X1 \ddin[7]$_DFFE_PN0P_  (
  .D(_019_),
  .RN(rst),
  .CK(clk),
  .Q(\ddin[8] ),
  .QN(_063_)
);

DFFR_X1 dgo$_DFFE_PN0P_ (
  .D(_008_),
  .RN(rst),
  .CK(clk),
  .Q(dgo),
  .QN(_074_)
);

DFFR_X1 douten$_DFFE_PN0P_ (
  .D(_006_),
  .RN(rst),
  .CK(clk),
  .Q(douten),
  .QN(_076_)
);

DFFR_X1 go$_DFFE_PN0P_ (
  .D(_007_),
  .RN(rst),
  .CK(clk),
  .Q(go),
  .QN(_075_)
);

DFFR_X1 \sample_cnt[0]$_DFFE_PN0P_  (
  .D(_000_),
  .RN(rst),
  .CK(clk),
  .Q(\sample_cnt[0] ),
  .QN(_082_)
);

DFFR_X1 \sample_cnt[1]$_DFFE_PN0P_  (
  .D(_001_),
  .RN(rst),
  .CK(clk),
  .Q(\sample_cnt[1] ),
  .QN(_081_)
);

DFFR_X1 \sample_cnt[2]$_DFFE_PN0P_  (
  .D(_002_),
  .RN(rst),
  .CK(clk),
  .Q(\sample_cnt[2] ),
  .QN(_080_)
);

DFFR_X1 \sample_cnt[3]$_DFFE_PN0P_  (
  .D(_003_),
  .RN(rst),
  .CK(clk),
  .Q(\sample_cnt[3] ),
  .QN(_079_)
);

DFFR_X1 \sample_cnt[4]$_DFFE_PN0P_  (
  .D(_004_),
  .RN(rst),
  .CK(clk),
  .Q(\sample_cnt[4] ),
  .QN(_078_)
);

DFFR_X1 \sample_cnt[5]$_DFFE_PN0P_  (
  .D(_005_),
  .RN(rst),
  .CK(clk),
  .Q(\sample_cnt[5] ),
  .QN(_077_)
);
endmodule //$paramod$849c8591669cf197b80ef99050b300773b555aae\dct

module \$paramod$849c8591669cf197b80ef99050b300773b555aae\fdct (input clk, input ena,
 input rst, input dstrb, input [7:0] din, output [11:0] dout, output douten);
wire doe;
wire \res00[0] ;
wire \res00[10] ;
wire \res00[11] ;
wire \res00[1] ;
wire \res00[2] ;
wire \res00[3] ;
wire \res00[4] ;
wire \res00[5] ;
wire \res00[6] ;
wire \res00[7] ;
wire \res00[8] ;
wire \res00[9] ;
wire \res01[0] ;
wire \res01[10] ;
wire \res01[11] ;
wire \res01[1] ;
wire \res01[2] ;
wire \res01[3] ;
wire \res01[4] ;
wire \res01[5] ;
wire \res01[6] ;
wire \res01[7] ;
wire \res01[8] ;
wire \res01[9] ;
wire \res02[0] ;
wire \res02[10] ;
wire \res02[11] ;
wire \res02[1] ;
wire \res02[2] ;
wire \res02[3] ;
wire \res02[4] ;
wire \res02[5] ;
wire \res02[6] ;
wire \res02[7] ;
wire \res02[8] ;
wire \res02[9] ;
wire \res03[0] ;
wire \res03[10] ;
wire \res03[11] ;
wire \res03[1] ;
wire \res03[2] ;
wire \res03[3] ;
wire \res03[4] ;
wire \res03[5] ;
wire \res03[6] ;
wire \res03[7] ;
wire \res03[8] ;
wire \res03[9] ;
wire \res04[0] ;
wire \res04[10] ;
wire \res04[11] ;
wire \res04[1] ;
wire \res04[2] ;
wire \res04[3] ;
wire \res04[4] ;
wire \res04[5] ;
wire \res04[6] ;
wire \res04[7] ;
wire \res04[8] ;
wire \res04[9] ;
wire \res05[0] ;
wire \res05[10] ;
wire \res05[11] ;
wire \res05[1] ;
wire \res05[2] ;
wire \res05[3] ;
wire \res05[4] ;
wire \res05[5] ;
wire \res05[6] ;
wire \res05[7] ;
wire \res05[8] ;
wire \res05[9] ;
wire \res06[0] ;
wire \res06[10] ;
wire \res06[11] ;
wire \res06[1] ;
wire \res06[2] ;
wire \res06[3] ;
wire \res06[4] ;
wire \res06[5] ;
wire \res06[6] ;
wire \res06[7] ;
wire \res06[8] ;
wire \res06[9] ;
wire \res07[0] ;
wire \res07[10] ;
wire \res07[11] ;
wire \res07[1] ;
wire \res07[2] ;
wire \res07[3] ;
wire \res07[4] ;
wire \res07[5] ;
wire \res07[6] ;
wire \res07[7] ;
wire \res07[8] ;
wire \res07[9] ;
wire \res10[0] ;
wire \res10[10] ;
wire \res10[11] ;
wire \res10[1] ;
wire \res10[2] ;
wire \res10[3] ;
wire \res10[4] ;
wire \res10[5] ;
wire \res10[6] ;
wire \res10[7] ;
wire \res10[8] ;
wire \res10[9] ;
wire \res11[0] ;
wire \res11[10] ;
wire \res11[11] ;
wire \res11[1] ;
wire \res11[2] ;
wire \res11[3] ;
wire \res11[4] ;
wire \res11[5] ;
wire \res11[6] ;
wire \res11[7] ;
wire \res11[8] ;
wire \res11[9] ;
wire \res12[0] ;
wire \res12[10] ;
wire \res12[11] ;
wire \res12[1] ;
wire \res12[2] ;
wire \res12[3] ;
wire \res12[4] ;
wire \res12[5] ;
wire \res12[6] ;
wire \res12[7] ;
wire \res12[8] ;
wire \res12[9] ;
wire \res13[0] ;
wire \res13[10] ;
wire \res13[11] ;
wire \res13[1] ;
wire \res13[2] ;
wire \res13[3] ;
wire \res13[4] ;
wire \res13[5] ;
wire \res13[6] ;
wire \res13[7] ;
wire \res13[8] ;
wire \res13[9] ;
wire \res14[0] ;
wire \res14[10] ;
wire \res14[11] ;
wire \res14[1] ;
wire \res14[2] ;
wire \res14[3] ;
wire \res14[4] ;
wire \res14[5] ;
wire \res14[6] ;
wire \res14[7] ;
wire \res14[8] ;
wire \res14[9] ;
wire \res15[0] ;
wire \res15[10] ;
wire \res15[11] ;
wire \res15[1] ;
wire \res15[2] ;
wire \res15[3] ;
wire \res15[4] ;
wire \res15[5] ;
wire \res15[6] ;
wire \res15[7] ;
wire \res15[8] ;
wire \res15[9] ;
wire \res16[0] ;
wire \res16[10] ;
wire \res16[11] ;
wire \res16[1] ;
wire \res16[2] ;
wire \res16[3] ;
wire \res16[4] ;
wire \res16[5] ;
wire \res16[6] ;
wire \res16[7] ;
wire \res16[8] ;
wire \res16[9] ;
wire \res17[0] ;
wire \res17[10] ;
wire \res17[11] ;
wire \res17[1] ;
wire \res17[2] ;
wire \res17[3] ;
wire \res17[4] ;
wire \res17[5] ;
wire \res17[6] ;
wire \res17[7] ;
wire \res17[8] ;
wire \res17[9] ;
wire \res20[0] ;
wire \res20[10] ;
wire \res20[11] ;
wire \res20[1] ;
wire \res20[2] ;
wire \res20[3] ;
wire \res20[4] ;
wire \res20[5] ;
wire \res20[6] ;
wire \res20[7] ;
wire \res20[8] ;
wire \res20[9] ;
wire \res21[0] ;
wire \res21[10] ;
wire \res21[11] ;
wire \res21[1] ;
wire \res21[2] ;
wire \res21[3] ;
wire \res21[4] ;
wire \res21[5] ;
wire \res21[6] ;
wire \res21[7] ;
wire \res21[8] ;
wire \res21[9] ;
wire \res22[0] ;
wire \res22[10] ;
wire \res22[11] ;
wire \res22[1] ;
wire \res22[2] ;
wire \res22[3] ;
wire \res22[4] ;
wire \res22[5] ;
wire \res22[6] ;
wire \res22[7] ;
wire \res22[8] ;
wire \res22[9] ;
wire \res23[0] ;
wire \res23[10] ;
wire \res23[11] ;
wire \res23[1] ;
wire \res23[2] ;
wire \res23[3] ;
wire \res23[4] ;
wire \res23[5] ;
wire \res23[6] ;
wire \res23[7] ;
wire \res23[8] ;
wire \res23[9] ;
wire \res24[0] ;
wire \res24[10] ;
wire \res24[11] ;
wire \res24[1] ;
wire \res24[2] ;
wire \res24[3] ;
wire \res24[4] ;
wire \res24[5] ;
wire \res24[6] ;
wire \res24[7] ;
wire \res24[8] ;
wire \res24[9] ;
wire \res25[0] ;
wire \res25[10] ;
wire \res25[11] ;
wire \res25[1] ;
wire \res25[2] ;
wire \res25[3] ;
wire \res25[4] ;
wire \res25[5] ;
wire \res25[6] ;
wire \res25[7] ;
wire \res25[8] ;
wire \res25[9] ;
wire \res26[0] ;
wire \res26[10] ;
wire \res26[11] ;
wire \res26[1] ;
wire \res26[2] ;
wire \res26[3] ;
wire \res26[4] ;
wire \res26[5] ;
wire \res26[6] ;
wire \res26[7] ;
wire \res26[8] ;
wire \res26[9] ;
wire \res27[0] ;
wire \res27[10] ;
wire \res27[11] ;
wire \res27[1] ;
wire \res27[2] ;
wire \res27[3] ;
wire \res27[4] ;
wire \res27[5] ;
wire \res27[6] ;
wire \res27[7] ;
wire \res27[8] ;
wire \res27[9] ;
wire \res30[0] ;
wire \res30[10] ;
wire \res30[11] ;
wire \res30[1] ;
wire \res30[2] ;
wire \res30[3] ;
wire \res30[4] ;
wire \res30[5] ;
wire \res30[6] ;
wire \res30[7] ;
wire \res30[8] ;
wire \res30[9] ;
wire \res31[0] ;
wire \res31[10] ;
wire \res31[11] ;
wire \res31[1] ;
wire \res31[2] ;
wire \res31[3] ;
wire \res31[4] ;
wire \res31[5] ;
wire \res31[6] ;
wire \res31[7] ;
wire \res31[8] ;
wire \res31[9] ;
wire \res32[0] ;
wire \res32[10] ;
wire \res32[11] ;
wire \res32[1] ;
wire \res32[2] ;
wire \res32[3] ;
wire \res32[4] ;
wire \res32[5] ;
wire \res32[6] ;
wire \res32[7] ;
wire \res32[8] ;
wire \res32[9] ;
wire \res33[0] ;
wire \res33[10] ;
wire \res33[11] ;
wire \res33[1] ;
wire \res33[2] ;
wire \res33[3] ;
wire \res33[4] ;
wire \res33[5] ;
wire \res33[6] ;
wire \res33[7] ;
wire \res33[8] ;
wire \res33[9] ;
wire \res34[0] ;
wire \res34[10] ;
wire \res34[11] ;
wire \res34[1] ;
wire \res34[2] ;
wire \res34[3] ;
wire \res34[4] ;
wire \res34[5] ;
wire \res34[6] ;
wire \res34[7] ;
wire \res34[8] ;
wire \res34[9] ;
wire \res35[0] ;
wire \res35[10] ;
wire \res35[11] ;
wire \res35[1] ;
wire \res35[2] ;
wire \res35[3] ;
wire \res35[4] ;
wire \res35[5] ;
wire \res35[6] ;
wire \res35[7] ;
wire \res35[8] ;
wire \res35[9] ;
wire \res36[0] ;
wire \res36[10] ;
wire \res36[11] ;
wire \res36[1] ;
wire \res36[2] ;
wire \res36[3] ;
wire \res36[4] ;
wire \res36[5] ;
wire \res36[6] ;
wire \res36[7] ;
wire \res36[8] ;
wire \res36[9] ;
wire \res37[0] ;
wire \res37[10] ;
wire \res37[11] ;
wire \res37[1] ;
wire \res37[2] ;
wire \res37[3] ;
wire \res37[4] ;
wire \res37[5] ;
wire \res37[6] ;
wire \res37[7] ;
wire \res37[8] ;
wire \res37[9] ;
wire \res40[0] ;
wire \res40[10] ;
wire \res40[11] ;
wire \res40[1] ;
wire \res40[2] ;
wire \res40[3] ;
wire \res40[4] ;
wire \res40[5] ;
wire \res40[6] ;
wire \res40[7] ;
wire \res40[8] ;
wire \res40[9] ;
wire \res41[0] ;
wire \res41[10] ;
wire \res41[11] ;
wire \res41[1] ;
wire \res41[2] ;
wire \res41[3] ;
wire \res41[4] ;
wire \res41[5] ;
wire \res41[6] ;
wire \res41[7] ;
wire \res41[8] ;
wire \res41[9] ;
wire \res42[0] ;
wire \res42[10] ;
wire \res42[11] ;
wire \res42[1] ;
wire \res42[2] ;
wire \res42[3] ;
wire \res42[4] ;
wire \res42[5] ;
wire \res42[6] ;
wire \res42[7] ;
wire \res42[8] ;
wire \res42[9] ;
wire \res43[0] ;
wire \res43[10] ;
wire \res43[11] ;
wire \res43[1] ;
wire \res43[2] ;
wire \res43[3] ;
wire \res43[4] ;
wire \res43[5] ;
wire \res43[6] ;
wire \res43[7] ;
wire \res43[8] ;
wire \res43[9] ;
wire \res44[0] ;
wire \res44[10] ;
wire \res44[11] ;
wire \res44[1] ;
wire \res44[2] ;
wire \res44[3] ;
wire \res44[4] ;
wire \res44[5] ;
wire \res44[6] ;
wire \res44[7] ;
wire \res44[8] ;
wire \res44[9] ;
wire \res45[0] ;
wire \res45[10] ;
wire \res45[11] ;
wire \res45[1] ;
wire \res45[2] ;
wire \res45[3] ;
wire \res45[4] ;
wire \res45[5] ;
wire \res45[6] ;
wire \res45[7] ;
wire \res45[8] ;
wire \res45[9] ;
wire \res46[0] ;
wire \res46[10] ;
wire \res46[11] ;
wire \res46[1] ;
wire \res46[2] ;
wire \res46[3] ;
wire \res46[4] ;
wire \res46[5] ;
wire \res46[6] ;
wire \res46[7] ;
wire \res46[8] ;
wire \res46[9] ;
wire \res47[0] ;
wire \res47[10] ;
wire \res47[11] ;
wire \res47[1] ;
wire \res47[2] ;
wire \res47[3] ;
wire \res47[4] ;
wire \res47[5] ;
wire \res47[6] ;
wire \res47[7] ;
wire \res47[8] ;
wire \res47[9] ;
wire \res50[0] ;
wire \res50[10] ;
wire \res50[11] ;
wire \res50[1] ;
wire \res50[2] ;
wire \res50[3] ;
wire \res50[4] ;
wire \res50[5] ;
wire \res50[6] ;
wire \res50[7] ;
wire \res50[8] ;
wire \res50[9] ;
wire \res51[0] ;
wire \res51[10] ;
wire \res51[11] ;
wire \res51[1] ;
wire \res51[2] ;
wire \res51[3] ;
wire \res51[4] ;
wire \res51[5] ;
wire \res51[6] ;
wire \res51[7] ;
wire \res51[8] ;
wire \res51[9] ;
wire \res52[0] ;
wire \res52[10] ;
wire \res52[11] ;
wire \res52[1] ;
wire \res52[2] ;
wire \res52[3] ;
wire \res52[4] ;
wire \res52[5] ;
wire \res52[6] ;
wire \res52[7] ;
wire \res52[8] ;
wire \res52[9] ;
wire \res53[0] ;
wire \res53[10] ;
wire \res53[11] ;
wire \res53[1] ;
wire \res53[2] ;
wire \res53[3] ;
wire \res53[4] ;
wire \res53[5] ;
wire \res53[6] ;
wire \res53[7] ;
wire \res53[8] ;
wire \res53[9] ;
wire \res54[0] ;
wire \res54[10] ;
wire \res54[11] ;
wire \res54[1] ;
wire \res54[2] ;
wire \res54[3] ;
wire \res54[4] ;
wire \res54[5] ;
wire \res54[6] ;
wire \res54[7] ;
wire \res54[8] ;
wire \res54[9] ;
wire \res55[0] ;
wire \res55[10] ;
wire \res55[11] ;
wire \res55[1] ;
wire \res55[2] ;
wire \res55[3] ;
wire \res55[4] ;
wire \res55[5] ;
wire \res55[6] ;
wire \res55[7] ;
wire \res55[8] ;
wire \res55[9] ;
wire \res56[0] ;
wire \res56[10] ;
wire \res56[11] ;
wire \res56[1] ;
wire \res56[2] ;
wire \res56[3] ;
wire \res56[4] ;
wire \res56[5] ;
wire \res56[6] ;
wire \res56[7] ;
wire \res56[8] ;
wire \res56[9] ;
wire \res57[0] ;
wire \res57[10] ;
wire \res57[11] ;
wire \res57[1] ;
wire \res57[2] ;
wire \res57[3] ;
wire \res57[4] ;
wire \res57[5] ;
wire \res57[6] ;
wire \res57[7] ;
wire \res57[8] ;
wire \res57[9] ;
wire \res60[0] ;
wire \res60[10] ;
wire \res60[11] ;
wire \res60[1] ;
wire \res60[2] ;
wire \res60[3] ;
wire \res60[4] ;
wire \res60[5] ;
wire \res60[6] ;
wire \res60[7] ;
wire \res60[8] ;
wire \res60[9] ;
wire \res61[0] ;
wire \res61[10] ;
wire \res61[11] ;
wire \res61[1] ;
wire \res61[2] ;
wire \res61[3] ;
wire \res61[4] ;
wire \res61[5] ;
wire \res61[6] ;
wire \res61[7] ;
wire \res61[8] ;
wire \res61[9] ;
wire \res62[0] ;
wire \res62[10] ;
wire \res62[11] ;
wire \res62[1] ;
wire \res62[2] ;
wire \res62[3] ;
wire \res62[4] ;
wire \res62[5] ;
wire \res62[6] ;
wire \res62[7] ;
wire \res62[8] ;
wire \res62[9] ;
wire \res63[0] ;
wire \res63[10] ;
wire \res63[11] ;
wire \res63[1] ;
wire \res63[2] ;
wire \res63[3] ;
wire \res63[4] ;
wire \res63[5] ;
wire \res63[6] ;
wire \res63[7] ;
wire \res63[8] ;
wire \res63[9] ;
wire \res64[0] ;
wire \res64[10] ;
wire \res64[11] ;
wire \res64[1] ;
wire \res64[2] ;
wire \res64[3] ;
wire \res64[4] ;
wire \res64[5] ;
wire \res64[6] ;
wire \res64[7] ;
wire \res64[8] ;
wire \res64[9] ;
wire \res65[0] ;
wire \res65[10] ;
wire \res65[11] ;
wire \res65[1] ;
wire \res65[2] ;
wire \res65[3] ;
wire \res65[4] ;
wire \res65[5] ;
wire \res65[6] ;
wire \res65[7] ;
wire \res65[8] ;
wire \res65[9] ;
wire \res66[0] ;
wire \res66[10] ;
wire \res66[11] ;
wire \res66[1] ;
wire \res66[2] ;
wire \res66[3] ;
wire \res66[4] ;
wire \res66[5] ;
wire \res66[6] ;
wire \res66[7] ;
wire \res66[8] ;
wire \res66[9] ;
wire \res67[0] ;
wire \res67[10] ;
wire \res67[11] ;
wire \res67[1] ;
wire \res67[2] ;
wire \res67[3] ;
wire \res67[4] ;
wire \res67[5] ;
wire \res67[6] ;
wire \res67[7] ;
wire \res67[8] ;
wire \res67[9] ;
wire \res70[0] ;
wire \res70[10] ;
wire \res70[11] ;
wire \res70[1] ;
wire \res70[2] ;
wire \res70[3] ;
wire \res70[4] ;
wire \res70[5] ;
wire \res70[6] ;
wire \res70[7] ;
wire \res70[8] ;
wire \res70[9] ;
wire \res71[0] ;
wire \res71[10] ;
wire \res71[11] ;
wire \res71[1] ;
wire \res71[2] ;
wire \res71[3] ;
wire \res71[4] ;
wire \res71[5] ;
wire \res71[6] ;
wire \res71[7] ;
wire \res71[8] ;
wire \res71[9] ;
wire \res72[0] ;
wire \res72[10] ;
wire \res72[11] ;
wire \res72[1] ;
wire \res72[2] ;
wire \res72[3] ;
wire \res72[4] ;
wire \res72[5] ;
wire \res72[6] ;
wire \res72[7] ;
wire \res72[8] ;
wire \res72[9] ;
wire \res73[0] ;
wire \res73[10] ;
wire \res73[11] ;
wire \res73[1] ;
wire \res73[2] ;
wire \res73[3] ;
wire \res73[4] ;
wire \res73[5] ;
wire \res73[6] ;
wire \res73[7] ;
wire \res73[8] ;
wire \res73[9] ;
wire \res74[0] ;
wire \res74[10] ;
wire \res74[11] ;
wire \res74[1] ;
wire \res74[2] ;
wire \res74[3] ;
wire \res74[4] ;
wire \res74[5] ;
wire \res74[6] ;
wire \res74[7] ;
wire \res74[8] ;
wire \res74[9] ;
wire \res75[0] ;
wire \res75[10] ;
wire \res75[11] ;
wire \res75[1] ;
wire \res75[2] ;
wire \res75[3] ;
wire \res75[4] ;
wire \res75[5] ;
wire \res75[6] ;
wire \res75[7] ;
wire \res75[8] ;
wire \res75[9] ;
wire \res76[0] ;
wire \res76[10] ;
wire \res76[11] ;
wire \res76[1] ;
wire \res76[2] ;
wire \res76[3] ;
wire \res76[4] ;
wire \res76[5] ;
wire \res76[6] ;
wire \res76[7] ;
wire \res76[8] ;
wire \res76[9] ;
wire \res77[0] ;
wire \res77[10] ;
wire \res77[11] ;
wire \res77[1] ;
wire \res77[2] ;
wire \res77[3] ;
wire \res77[4] ;
wire \res77[5] ;
wire \res77[6] ;
wire \res77[7] ;
wire \res77[8] ;
wire \res77[9] ;

\$paramod$849c8591669cf197b80ef99050b300773b555aae\dct  dct_mod (
  .clk(clk),
  .ena(ena),
  .rst(rst),
  .dstrb(dstrb),
  .din(din),
  .dout_00({\res00[11] , \res00[10] , \res00[9] , \res00[8] , \res00[7] , \res00[6] , \res00[5] , \res00[4] , \res00[3] , \res00[2] , \res00[1] , \res00[0] }),
  .dout_01({\res01[11] , \res01[10] , \res01[9] , \res01[8] , \res01[7] , \res01[6] , \res01[5] , \res01[4] , \res01[3] , \res01[2] , \res01[1] , \res01[0] }),
  .dout_02({\res02[11] , \res02[10] , \res02[9] , \res02[8] , \res02[7] , \res02[6] , \res02[5] , \res02[4] , \res02[3] , \res02[2] , \res02[1] , \res02[0] }),
  .dout_03({\res03[11] , \res03[10] , \res03[9] , \res03[8] , \res03[7] , \res03[6] , \res03[5] , \res03[4] , \res03[3] , \res03[2] , \res03[1] , \res03[0] }),
  .dout_04({\res04[11] , \res04[10] , \res04[9] , \res04[8] , \res04[7] , \res04[6] , \res04[5] , \res04[4] , \res04[3] , \res04[2] , \res04[1] , \res04[0] }),
  .dout_05({\res05[11] , \res05[10] , \res05[9] , \res05[8] , \res05[7] , \res05[6] , \res05[5] , \res05[4] , \res05[3] , \res05[2] , \res05[1] , \res05[0] }),
  .dout_06({\res06[11] , \res06[10] , \res06[9] , \res06[8] , \res06[7] , \res06[6] , \res06[5] , \res06[4] , \res06[3] , \res06[2] , \res06[1] , \res06[0] }),
  .dout_07({\res07[11] , \res07[10] , \res07[9] , \res07[8] , \res07[7] , \res07[6] , \res07[5] , \res07[4] , \res07[3] , \res07[2] , \res07[1] , \res07[0] }),
  .dout_10({\res10[11] , \res10[10] , \res10[9] , \res10[8] , \res10[7] , \res10[6] , \res10[5] , \res10[4] , \res10[3] , \res10[2] , \res10[1] , \res10[0] }),
  .dout_11({\res11[11] , \res11[10] , \res11[9] , \res11[8] , \res11[7] , \res11[6] , \res11[5] , \res11[4] , \res11[3] , \res11[2] , \res11[1] , \res11[0] }),
  .dout_12({\res12[11] , \res12[10] , \res12[9] , \res12[8] , \res12[7] , \res12[6] , \res12[5] , \res12[4] , \res12[3] , \res12[2] , \res12[1] , \res12[0] }),
  .dout_13({\res13[11] , \res13[10] , \res13[9] , \res13[8] , \res13[7] , \res13[6] , \res13[5] , \res13[4] , \res13[3] , \res13[2] , \res13[1] , \res13[0] }),
  .dout_14({\res14[11] , \res14[10] , \res14[9] , \res14[8] , \res14[7] , \res14[6] , \res14[5] , \res14[4] , \res14[3] , \res14[2] , \res14[1] , \res14[0] }),
  .dout_15({\res15[11] , \res15[10] , \res15[9] , \res15[8] , \res15[7] , \res15[6] , \res15[5] , \res15[4] , \res15[3] , \res15[2] , \res15[1] , \res15[0] }),
  .dout_16({\res16[11] , \res16[10] , \res16[9] , \res16[8] , \res16[7] , \res16[6] , \res16[5] , \res16[4] , \res16[3] , \res16[2] , \res16[1] , \res16[0] }),
  .dout_17({\res17[11] , \res17[10] , \res17[9] , \res17[8] , \res17[7] , \res17[6] , \res17[5] , \res17[4] , \res17[3] , \res17[2] , \res17[1] , \res17[0] }),
  .dout_20({\res20[11] , \res20[10] , \res20[9] , \res20[8] , \res20[7] , \res20[6] , \res20[5] , \res20[4] , \res20[3] , \res20[2] , \res20[1] , \res20[0] }),
  .dout_21({\res21[11] , \res21[10] , \res21[9] , \res21[8] , \res21[7] , \res21[6] , \res21[5] , \res21[4] , \res21[3] , \res21[2] , \res21[1] , \res21[0] }),
  .dout_22({\res22[11] , \res22[10] , \res22[9] , \res22[8] , \res22[7] , \res22[6] , \res22[5] , \res22[4] , \res22[3] , \res22[2] , \res22[1] , \res22[0] }),
  .dout_23({\res23[11] , \res23[10] , \res23[9] , \res23[8] , \res23[7] , \res23[6] , \res23[5] , \res23[4] , \res23[3] , \res23[2] , \res23[1] , \res23[0] }),
  .dout_24({\res24[11] , \res24[10] , \res24[9] , \res24[8] , \res24[7] , \res24[6] , \res24[5] , \res24[4] , \res24[3] , \res24[2] , \res24[1] , \res24[0] }),
  .dout_25({\res25[11] , \res25[10] , \res25[9] , \res25[8] , \res25[7] , \res25[6] , \res25[5] , \res25[4] , \res25[3] , \res25[2] , \res25[1] , \res25[0] }),
  .dout_26({\res26[11] , \res26[10] , \res26[9] , \res26[8] , \res26[7] , \res26[6] , \res26[5] , \res26[4] , \res26[3] , \res26[2] , \res26[1] , \res26[0] }),
  .dout_27({\res27[11] , \res27[10] , \res27[9] , \res27[8] , \res27[7] , \res27[6] , \res27[5] , \res27[4] , \res27[3] , \res27[2] , \res27[1] , \res27[0] }),
  .dout_30({\res30[11] , \res30[10] , \res30[9] , \res30[8] , \res30[7] , \res30[6] , \res30[5] , \res30[4] , \res30[3] , \res30[2] , \res30[1] , \res30[0] }),
  .dout_31({\res31[11] , \res31[10] , \res31[9] , \res31[8] , \res31[7] , \res31[6] , \res31[5] , \res31[4] , \res31[3] , \res31[2] , \res31[1] , \res31[0] }),
  .dout_32({\res32[11] , \res32[10] , \res32[9] , \res32[8] , \res32[7] , \res32[6] , \res32[5] , \res32[4] , \res32[3] , \res32[2] , \res32[1] , \res32[0] }),
  .dout_33({\res33[11] , \res33[10] , \res33[9] , \res33[8] , \res33[7] , \res33[6] , \res33[5] , \res33[4] , \res33[3] , \res33[2] , \res33[1] , \res33[0] }),
  .dout_34({\res34[11] , \res34[10] , \res34[9] , \res34[8] , \res34[7] , \res34[6] , \res34[5] , \res34[4] , \res34[3] , \res34[2] , \res34[1] , \res34[0] }),
  .dout_35({\res35[11] , \res35[10] , \res35[9] , \res35[8] , \res35[7] , \res35[6] , \res35[5] , \res35[4] , \res35[3] , \res35[2] , \res35[1] , \res35[0] }),
  .dout_36({\res36[11] , \res36[10] , \res36[9] , \res36[8] , \res36[7] , \res36[6] , \res36[5] , \res36[4] , \res36[3] , \res36[2] , \res36[1] , \res36[0] }),
  .dout_37({\res37[11] , \res37[10] , \res37[9] , \res37[8] , \res37[7] , \res37[6] , \res37[5] , \res37[4] , \res37[3] , \res37[2] , \res37[1] , \res37[0] }),
  .dout_40({\res40[11] , \res40[10] , \res40[9] , \res40[8] , \res40[7] , \res40[6] , \res40[5] , \res40[4] , \res40[3] , \res40[2] , \res40[1] , \res40[0] }),
  .dout_41({\res41[11] , \res41[10] , \res41[9] , \res41[8] , \res41[7] , \res41[6] , \res41[5] , \res41[4] , \res41[3] , \res41[2] , \res41[1] , \res41[0] }),
  .dout_42({\res42[11] , \res42[10] , \res42[9] , \res42[8] , \res42[7] , \res42[6] , \res42[5] , \res42[4] , \res42[3] , \res42[2] , \res42[1] , \res42[0] }),
  .dout_43({\res43[11] , \res43[10] , \res43[9] , \res43[8] , \res43[7] , \res43[6] , \res43[5] , \res43[4] , \res43[3] , \res43[2] , \res43[1] , \res43[0] }),
  .dout_44({\res44[11] , \res44[10] , \res44[9] , \res44[8] , \res44[7] , \res44[6] , \res44[5] , \res44[4] , \res44[3] , \res44[2] , \res44[1] , \res44[0] }),
  .dout_45({\res45[11] , \res45[10] , \res45[9] , \res45[8] , \res45[7] , \res45[6] , \res45[5] , \res45[4] , \res45[3] , \res45[2] , \res45[1] , \res45[0] }),
  .dout_46({\res46[11] , \res46[10] , \res46[9] , \res46[8] , \res46[7] , \res46[6] , \res46[5] , \res46[4] , \res46[3] , \res46[2] , \res46[1] , \res46[0] }),
  .dout_47({\res47[11] , \res47[10] , \res47[9] , \res47[8] , \res47[7] , \res47[6] , \res47[5] , \res47[4] , \res47[3] , \res47[2] , \res47[1] , \res47[0] }),
  .dout_50({\res50[11] , \res50[10] , \res50[9] , \res50[8] , \res50[7] , \res50[6] , \res50[5] , \res50[4] , \res50[3] , \res50[2] , \res50[1] , \res50[0] }),
  .dout_51({\res51[11] , \res51[10] , \res51[9] , \res51[8] , \res51[7] , \res51[6] , \res51[5] , \res51[4] , \res51[3] , \res51[2] , \res51[1] , \res51[0] }),
  .dout_52({\res52[11] , \res52[10] , \res52[9] , \res52[8] , \res52[7] , \res52[6] , \res52[5] , \res52[4] , \res52[3] , \res52[2] , \res52[1] , \res52[0] }),
  .dout_53({\res53[11] , \res53[10] , \res53[9] , \res53[8] , \res53[7] , \res53[6] , \res53[5] , \res53[4] , \res53[3] , \res53[2] , \res53[1] , \res53[0] }),
  .dout_54({\res54[11] , \res54[10] , \res54[9] , \res54[8] , \res54[7] , \res54[6] , \res54[5] , \res54[4] , \res54[3] , \res54[2] , \res54[1] , \res54[0] }),
  .dout_55({\res55[11] , \res55[10] , \res55[9] , \res55[8] , \res55[7] , \res55[6] , \res55[5] , \res55[4] , \res55[3] , \res55[2] , \res55[1] , \res55[0] }),
  .dout_56({\res56[11] , \res56[10] , \res56[9] , \res56[8] , \res56[7] , \res56[6] , \res56[5] , \res56[4] , \res56[3] , \res56[2] , \res56[1] , \res56[0] }),
  .dout_57({\res57[11] , \res57[10] , \res57[9] , \res57[8] , \res57[7] , \res57[6] , \res57[5] , \res57[4] , \res57[3] , \res57[2] , \res57[1] , \res57[0] }),
  .dout_60({\res60[11] , \res60[10] , \res60[9] , \res60[8] , \res60[7] , \res60[6] , \res60[5] , \res60[4] , \res60[3] , \res60[2] , \res60[1] , \res60[0] }),
  .dout_61({\res61[11] , \res61[10] , \res61[9] , \res61[8] , \res61[7] , \res61[6] , \res61[5] , \res61[4] , \res61[3] , \res61[2] , \res61[1] , \res61[0] }),
  .dout_62({\res62[11] , \res62[10] , \res62[9] , \res62[8] , \res62[7] , \res62[6] , \res62[5] , \res62[4] , \res62[3] , \res62[2] , \res62[1] , \res62[0] }),
  .dout_63({\res63[11] , \res63[10] , \res63[9] , \res63[8] , \res63[7] , \res63[6] , \res63[5] , \res63[4] , \res63[3] , \res63[2] , \res63[1] , \res63[0] }),
  .dout_64({\res64[11] , \res64[10] , \res64[9] , \res64[8] , \res64[7] , \res64[6] , \res64[5] , \res64[4] , \res64[3] , \res64[2] , \res64[1] , \res64[0] }),
  .dout_65({\res65[11] , \res65[10] , \res65[9] , \res65[8] , \res65[7] , \res65[6] , \res65[5] , \res65[4] , \res65[3] , \res65[2] , \res65[1] , \res65[0] }),
  .dout_66({\res66[11] , \res66[10] , \res66[9] , \res66[8] , \res66[7] , \res66[6] , \res66[5] , \res66[4] , \res66[3] , \res66[2] , \res66[1] , \res66[0] }),
  .dout_67({\res67[11] , \res67[10] , \res67[9] , \res67[8] , \res67[7] , \res67[6] , \res67[5] , \res67[4] , \res67[3] , \res67[2] , \res67[1] , \res67[0] }),
  .dout_70({\res70[11] , \res70[10] , \res70[9] , \res70[8] , \res70[7] , \res70[6] , \res70[5] , \res70[4] , \res70[3] , \res70[2] , \res70[1] , \res70[0] }),
  .dout_71({\res71[11] , \res71[10] , \res71[9] , \res71[8] , \res71[7] , \res71[6] , \res71[5] , \res71[4] , \res71[3] , \res71[2] , \res71[1] , \res71[0] }),
  .dout_72({\res72[11] , \res72[10] , \res72[9] , \res72[8] , \res72[7] , \res72[6] , \res72[5] , \res72[4] , \res72[3] , \res72[2] , \res72[1] , \res72[0] }),
  .dout_73({\res73[11] , \res73[10] , \res73[9] , \res73[8] , \res73[7] , \res73[6] , \res73[5] , \res73[4] , \res73[3] , \res73[2] , \res73[1] , \res73[0] }),
  .dout_74({\res74[11] , \res74[10] , \res74[9] , \res74[8] , \res74[7] , \res74[6] , \res74[5] , \res74[4] , \res74[3] , \res74[2] , \res74[1] , \res74[0] }),
  .dout_75({\res75[11] , \res75[10] , \res75[9] , \res75[8] , \res75[7] , \res75[6] , \res75[5] , \res75[4] , \res75[3] , \res75[2] , \res75[1] , \res75[0] }),
  .dout_76({\res76[11] , \res76[10] , \res76[9] , \res76[8] , \res76[7] , \res76[6] , \res76[5] , \res76[4] , \res76[3] , \res76[2] , \res76[1] , \res76[0] }),
  .dout_77({\res77[11] , \res77[10] , \res77[9] , \res77[8] , \res77[7] , \res77[6] , \res77[5] , \res77[4] , \res77[3] , \res77[2] , \res77[1] , \res77[0] }),
  .douten(doe)
);

zigzag zigzag_mod (
  .clk(clk),
  .ena(ena),
  .dstrb(doe),
  .din_00({\res00[11] , \res00[10] , \res00[9] , \res00[8] , \res00[7] , \res00[6] , \res00[5] , \res00[4] , \res00[3] , \res00[2] , \res00[1] , \res00[0] }),
  .din_01({\res01[11] , \res01[10] , \res01[9] , \res01[8] , \res01[7] , \res01[6] , \res01[5] , \res01[4] , \res01[3] , \res01[2] , \res01[1] , \res01[0] }),
  .din_02({\res02[11] , \res02[10] , \res02[9] , \res02[8] , \res02[7] , \res02[6] , \res02[5] , \res02[4] , \res02[3] , \res02[2] , \res02[1] , \res02[0] }),
  .din_03({\res03[11] , \res03[10] , \res03[9] , \res03[8] , \res03[7] , \res03[6] , \res03[5] , \res03[4] , \res03[3] , \res03[2] , \res03[1] , \res03[0] }),
  .din_04({\res04[11] , \res04[10] , \res04[9] , \res04[8] , \res04[7] , \res04[6] , \res04[5] , \res04[4] , \res04[3] , \res04[2] , \res04[1] , \res04[0] }),
  .din_05({\res05[11] , \res05[10] , \res05[9] , \res05[8] , \res05[7] , \res05[6] , \res05[5] , \res05[4] , \res05[3] , \res05[2] , \res05[1] , \res05[0] }),
  .din_06({\res06[11] , \res06[10] , \res06[9] , \res06[8] , \res06[7] , \res06[6] , \res06[5] , \res06[4] , \res06[3] , \res06[2] , \res06[1] , \res06[0] }),
  .din_07({\res07[11] , \res07[10] , \res07[9] , \res07[8] , \res07[7] , \res07[6] , \res07[5] , \res07[4] , \res07[3] , \res07[2] , \res07[1] , \res07[0] }),
  .din_10({\res10[11] , \res10[10] , \res10[9] , \res10[8] , \res10[7] , \res10[6] , \res10[5] , \res10[4] , \res10[3] , \res10[2] , \res10[1] , \res10[0] }),
  .din_11({\res11[11] , \res11[10] , \res11[9] , \res11[8] , \res11[7] , \res11[6] , \res11[5] , \res11[4] , \res11[3] , \res11[2] , \res11[1] , \res11[0] }),
  .din_12({\res12[11] , \res12[10] , \res12[9] , \res12[8] , \res12[7] , \res12[6] , \res12[5] , \res12[4] , \res12[3] , \res12[2] , \res12[1] , \res12[0] }),
  .din_13({\res13[11] , \res13[10] , \res13[9] , \res13[8] , \res13[7] , \res13[6] , \res13[5] , \res13[4] , \res13[3] , \res13[2] , \res13[1] , \res13[0] }),
  .din_14({\res14[11] , \res14[10] , \res14[9] , \res14[8] , \res14[7] , \res14[6] , \res14[5] , \res14[4] , \res14[3] , \res14[2] , \res14[1] , \res14[0] }),
  .din_15({\res15[11] , \res15[10] , \res15[9] , \res15[8] , \res15[7] , \res15[6] , \res15[5] , \res15[4] , \res15[3] , \res15[2] , \res15[1] , \res15[0] }),
  .din_16({\res16[11] , \res16[10] , \res16[9] , \res16[8] , \res16[7] , \res16[6] , \res16[5] , \res16[4] , \res16[3] , \res16[2] , \res16[1] , \res16[0] }),
  .din_17({\res17[11] , \res17[10] , \res17[9] , \res17[8] , \res17[7] , \res17[6] , \res17[5] , \res17[4] , \res17[3] , \res17[2] , \res17[1] , \res17[0] }),
  .din_20({\res20[11] , \res20[10] , \res20[9] , \res20[8] , \res20[7] , \res20[6] , \res20[5] , \res20[4] , \res20[3] , \res20[2] , \res20[1] , \res20[0] }),
  .din_21({\res21[11] , \res21[10] , \res21[9] , \res21[8] , \res21[7] , \res21[6] , \res21[5] , \res21[4] , \res21[3] , \res21[2] , \res21[1] , \res21[0] }),
  .din_22({\res22[11] , \res22[10] , \res22[9] , \res22[8] , \res22[7] , \res22[6] , \res22[5] , \res22[4] , \res22[3] , \res22[2] , \res22[1] , \res22[0] }),
  .din_23({\res23[11] , \res23[10] , \res23[9] , \res23[8] , \res23[7] , \res23[6] , \res23[5] , \res23[4] , \res23[3] , \res23[2] , \res23[1] , \res23[0] }),
  .din_24({\res24[11] , \res24[10] , \res24[9] , \res24[8] , \res24[7] , \res24[6] , \res24[5] , \res24[4] , \res24[3] , \res24[2] , \res24[1] , \res24[0] }),
  .din_25({\res25[11] , \res25[10] , \res25[9] , \res25[8] , \res25[7] , \res25[6] , \res25[5] , \res25[4] , \res25[3] , \res25[2] , \res25[1] , \res25[0] }),
  .din_26({\res26[11] , \res26[10] , \res26[9] , \res26[8] , \res26[7] , \res26[6] , \res26[5] , \res26[4] , \res26[3] , \res26[2] , \res26[1] , \res26[0] }),
  .din_27({\res27[11] , \res27[10] , \res27[9] , \res27[8] , \res27[7] , \res27[6] , \res27[5] , \res27[4] , \res27[3] , \res27[2] , \res27[1] , \res27[0] }),
  .din_30({\res30[11] , \res30[10] , \res30[9] , \res30[8] , \res30[7] , \res30[6] , \res30[5] , \res30[4] , \res30[3] , \res30[2] , \res30[1] , \res30[0] }),
  .din_31({\res31[11] , \res31[10] , \res31[9] , \res31[8] , \res31[7] , \res31[6] , \res31[5] , \res31[4] , \res31[3] , \res31[2] , \res31[1] , \res31[0] }),
  .din_32({\res32[11] , \res32[10] , \res32[9] , \res32[8] , \res32[7] , \res32[6] , \res32[5] , \res32[4] , \res32[3] , \res32[2] , \res32[1] , \res32[0] }),
  .din_33({\res33[11] , \res33[10] , \res33[9] , \res33[8] , \res33[7] , \res33[6] , \res33[5] , \res33[4] , \res33[3] , \res33[2] , \res33[1] , \res33[0] }),
  .din_34({\res34[11] , \res34[10] , \res34[9] , \res34[8] , \res34[7] , \res34[6] , \res34[5] , \res34[4] , \res34[3] , \res34[2] , \res34[1] , \res34[0] }),
  .din_35({\res35[11] , \res35[10] , \res35[9] , \res35[8] , \res35[7] , \res35[6] , \res35[5] , \res35[4] , \res35[3] , \res35[2] , \res35[1] , \res35[0] }),
  .din_36({\res36[11] , \res36[10] , \res36[9] , \res36[8] , \res36[7] , \res36[6] , \res36[5] , \res36[4] , \res36[3] , \res36[2] , \res36[1] , \res36[0] }),
  .din_37({\res37[11] , \res37[10] , \res37[9] , \res37[8] , \res37[7] , \res37[6] , \res37[5] , \res37[4] , \res37[3] , \res37[2] , \res37[1] , \res37[0] }),
  .din_40({\res40[11] , \res40[10] , \res40[9] , \res40[8] , \res40[7] , \res40[6] , \res40[5] , \res40[4] , \res40[3] , \res40[2] , \res40[1] , \res40[0] }),
  .din_41({\res41[11] , \res41[10] , \res41[9] , \res41[8] , \res41[7] , \res41[6] , \res41[5] , \res41[4] , \res41[3] , \res41[2] , \res41[1] , \res41[0] }),
  .din_42({\res42[11] , \res42[10] , \res42[9] , \res42[8] , \res42[7] , \res42[6] , \res42[5] , \res42[4] , \res42[3] , \res42[2] , \res42[1] , \res42[0] }),
  .din_43({\res43[11] , \res43[10] , \res43[9] , \res43[8] , \res43[7] , \res43[6] , \res43[5] , \res43[4] , \res43[3] , \res43[2] , \res43[1] , \res43[0] }),
  .din_44({\res44[11] , \res44[10] , \res44[9] , \res44[8] , \res44[7] , \res44[6] , \res44[5] , \res44[4] , \res44[3] , \res44[2] , \res44[1] , \res44[0] }),
  .din_45({\res45[11] , \res45[10] , \res45[9] , \res45[8] , \res45[7] , \res45[6] , \res45[5] , \res45[4] , \res45[3] , \res45[2] , \res45[1] , \res45[0] }),
  .din_46({\res46[11] , \res46[10] , \res46[9] , \res46[8] , \res46[7] , \res46[6] , \res46[5] , \res46[4] , \res46[3] , \res46[2] , \res46[1] , \res46[0] }),
  .din_47({\res47[11] , \res47[10] , \res47[9] , \res47[8] , \res47[7] , \res47[6] , \res47[5] , \res47[4] , \res47[3] , \res47[2] , \res47[1] , \res47[0] }),
  .din_50({\res50[11] , \res50[10] , \res50[9] , \res50[8] , \res50[7] , \res50[6] , \res50[5] , \res50[4] , \res50[3] , \res50[2] , \res50[1] , \res50[0] }),
  .din_51({\res51[11] , \res51[10] , \res51[9] , \res51[8] , \res51[7] , \res51[6] , \res51[5] , \res51[4] , \res51[3] , \res51[2] , \res51[1] , \res51[0] }),
  .din_52({\res52[11] , \res52[10] , \res52[9] , \res52[8] , \res52[7] , \res52[6] , \res52[5] , \res52[4] , \res52[3] , \res52[2] , \res52[1] , \res52[0] }),
  .din_53({\res53[11] , \res53[10] , \res53[9] , \res53[8] , \res53[7] , \res53[6] , \res53[5] , \res53[4] , \res53[3] , \res53[2] , \res53[1] , \res53[0] }),
  .din_54({\res54[11] , \res54[10] , \res54[9] , \res54[8] , \res54[7] , \res54[6] , \res54[5] , \res54[4] , \res54[3] , \res54[2] , \res54[1] , \res54[0] }),
  .din_55({\res55[11] , \res55[10] , \res55[9] , \res55[8] , \res55[7] , \res55[6] , \res55[5] , \res55[4] , \res55[3] , \res55[2] , \res55[1] , \res55[0] }),
  .din_56({\res56[11] , \res56[10] , \res56[9] , \res56[8] , \res56[7] , \res56[6] , \res56[5] , \res56[4] , \res56[3] , \res56[2] , \res56[1] , \res56[0] }),
  .din_57({\res57[11] , \res57[10] , \res57[9] , \res57[8] , \res57[7] , \res57[6] , \res57[5] , \res57[4] , \res57[3] , \res57[2] , \res57[1] , \res57[0] }),
  .din_60({\res60[11] , \res60[10] , \res60[9] , \res60[8] , \res60[7] , \res60[6] , \res60[5] , \res60[4] , \res60[3] , \res60[2] , \res60[1] , \res60[0] }),
  .din_61({\res61[11] , \res61[10] , \res61[9] , \res61[8] , \res61[7] , \res61[6] , \res61[5] , \res61[4] , \res61[3] , \res61[2] , \res61[1] , \res61[0] }),
  .din_62({\res62[11] , \res62[10] , \res62[9] , \res62[8] , \res62[7] , \res62[6] , \res62[5] , \res62[4] , \res62[3] , \res62[2] , \res62[1] , \res62[0] }),
  .din_63({\res63[11] , \res63[10] , \res63[9] , \res63[8] , \res63[7] , \res63[6] , \res63[5] , \res63[4] , \res63[3] , \res63[2] , \res63[1] , \res63[0] }),
  .din_64({\res64[11] , \res64[10] , \res64[9] , \res64[8] , \res64[7] , \res64[6] , \res64[5] , \res64[4] , \res64[3] , \res64[2] , \res64[1] , \res64[0] }),
  .din_65({\res65[11] , \res65[10] , \res65[9] , \res65[8] , \res65[7] , \res65[6] , \res65[5] , \res65[4] , \res65[3] , \res65[2] , \res65[1] , \res65[0] }),
  .din_66({\res66[11] , \res66[10] , \res66[9] , \res66[8] , \res66[7] , \res66[6] , \res66[5] , \res66[4] , \res66[3] , \res66[2] , \res66[1] , \res66[0] }),
  .din_67({\res67[11] , \res67[10] , \res67[9] , \res67[8] , \res67[7] , \res67[6] , \res67[5] , \res67[4] , \res67[3] , \res67[2] , \res67[1] , \res67[0] }),
  .din_70({\res70[11] , \res70[10] , \res70[9] , \res70[8] , \res70[7] , \res70[6] , \res70[5] , \res70[4] , \res70[3] , \res70[2] , \res70[1] , \res70[0] }),
  .din_71({\res71[11] , \res71[10] , \res71[9] , \res71[8] , \res71[7] , \res71[6] , \res71[5] , \res71[4] , \res71[3] , \res71[2] , \res71[1] , \res71[0] }),
  .din_72({\res72[11] , \res72[10] , \res72[9] , \res72[8] , \res72[7] , \res72[6] , \res72[5] , \res72[4] , \res72[3] , \res72[2] , \res72[1] , \res72[0] }),
  .din_73({\res73[11] , \res73[10] , \res73[9] , \res73[8] , \res73[7] , \res73[6] , \res73[5] , \res73[4] , \res73[3] , \res73[2] , \res73[1] , \res73[0] }),
  .din_74({\res74[11] , \res74[10] , \res74[9] , \res74[8] , \res74[7] , \res74[6] , \res74[5] , \res74[4] , \res74[3] , \res74[2] , \res74[1] , \res74[0] }),
  .din_75({\res75[11] , \res75[10] , \res75[9] , \res75[8] , \res75[7] , \res75[6] , \res75[5] , \res75[4] , \res75[3] , \res75[2] , \res75[1] , \res75[0] }),
  .din_76({\res76[11] , \res76[10] , \res76[9] , \res76[8] , \res76[7] , \res76[6] , \res76[5] , \res76[4] , \res76[3] , \res76[2] , \res76[1] , \res76[0] }),
  .din_77({\res77[11] , \res77[10] , \res77[9] , \res77[8] , \res77[7] , \res77[6] , \res77[5] , \res77[4] , \res77[3] , \res77[2] , \res77[1] , \res77[0] }),
  .dout(dout),
  .douten(douten)
);
endmodule //$paramod$849c8591669cf197b80ef99050b300773b555aae\fdct

module jpeg_encoder(input clk, input ena, input rst, input dstrb, input [7:0] din,
 input [7:0] qnt_val, output [5:0] qnt_cnt, output [3:0] size, output [3:0] rlen, output [11:0] amp,
 output douten);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire dc_diff_doe;
wire \dfdct_dout[0] ;
wire \dfdct_dout[10] ;
wire \dfdct_dout[11] ;
wire \dfdct_dout[1] ;
wire \dfdct_dout[2] ;
wire \dfdct_dout[3] ;
wire \dfdct_dout[4] ;
wire \dfdct_dout[5] ;
wire \dfdct_dout[6] ;
wire \dfdct_dout[7] ;
wire \dfdct_dout[8] ;
wire \dfdct_dout[9] ;
wire fdct_doe;
wire \fdct_dout[0] ;
wire \fdct_dout[10] ;
wire \fdct_dout[11] ;
wire \fdct_dout[1] ;
wire \fdct_dout[2] ;
wire \fdct_dout[3] ;
wire \fdct_dout[4] ;
wire \fdct_dout[5] ;
wire \fdct_dout[6] ;
wire \fdct_dout[7] ;
wire \fdct_dout[8] ;
wire \fdct_dout[9] ;
wire qnr_doe;
wire \qnr_dout[0] ;
wire \qnr_dout[10] ;
wire \qnr_dout[1] ;
wire \qnr_dout[2] ;
wire \qnr_dout[3] ;
wire \qnr_dout[4] ;
wire \qnr_dout[5] ;
wire \qnr_dout[6] ;
wire \qnr_dout[7] ;
wire \qnr_dout[8] ;
wire \qnr_dout[9] ;

BUF_X4 _56_ (
  .A(ena),
  .Z(_13_)
);

INV_X8 _57_ (
  .A(_13_),
  .ZN(_14_)
);

BUF_X32 _58_ (
  .A(_14_),
  .Z(_15_)
);

NAND2_X4 _59_ (
  .A1(_15_),
  .A2(\dfdct_dout[0] ),
  .ZN(_16_)
);

NAND2_X1 _60_ (
  .A1(\fdct_dout[0] ),
  .A2(_13_),
  .ZN(_17_)
);

NAND2_X4 _61_ (
  .A1(_16_),
  .A2(_17_),
  .ZN(_00_)
);

NAND2_X4 _62_ (
  .A1(_15_),
  .A2(\dfdct_dout[2] ),
  .ZN(_18_)
);

BUF_X8 _63_ (
  .A(_13_),
  .Z(_19_)
);

NAND2_X1 _64_ (
  .A1(_19_),
  .A2(\fdct_dout[2] ),
  .ZN(_20_)
);

NAND2_X2 _65_ (
  .A1(_18_),
  .A2(_20_),
  .ZN(_01_)
);

NAND2_X4 _66_ (
  .A1(_15_),
  .A2(\dfdct_dout[3] ),
  .ZN(_21_)
);

NAND2_X1 _67_ (
  .A1(_19_),
  .A2(\fdct_dout[3] ),
  .ZN(_22_)
);

NAND2_X2 _68_ (
  .A1(_21_),
  .A2(_22_),
  .ZN(_02_)
);

NAND2_X4 _69_ (
  .A1(_15_),
  .A2(\dfdct_dout[4] ),
  .ZN(_23_)
);

NAND2_X1 _70_ (
  .A1(_19_),
  .A2(\fdct_dout[4] ),
  .ZN(_24_)
);

NAND2_X2 _71_ (
  .A1(_23_),
  .A2(_24_),
  .ZN(_03_)
);

NAND2_X4 _72_ (
  .A1(_15_),
  .A2(\dfdct_dout[5] ),
  .ZN(_25_)
);

NAND2_X1 _73_ (
  .A1(_13_),
  .A2(\fdct_dout[5] ),
  .ZN(_26_)
);

NAND2_X4 _74_ (
  .A1(_25_),
  .A2(_26_),
  .ZN(_04_)
);

NAND2_X4 _75_ (
  .A1(_15_),
  .A2(\dfdct_dout[6] ),
  .ZN(_27_)
);

NAND2_X1 _76_ (
  .A1(_19_),
  .A2(\fdct_dout[6] ),
  .ZN(_28_)
);

NAND2_X2 _77_ (
  .A1(_27_),
  .A2(_28_),
  .ZN(_05_)
);

NAND2_X1 _78_ (
  .A1(_14_),
  .A2(\dfdct_dout[7] ),
  .ZN(_29_)
);

NAND2_X1 _79_ (
  .A1(_19_),
  .A2(\fdct_dout[7] ),
  .ZN(_30_)
);

NAND2_X1 _80_ (
  .A1(_29_),
  .A2(_30_),
  .ZN(_06_)
);

NAND2_X4 _81_ (
  .A1(_15_),
  .A2(\dfdct_dout[8] ),
  .ZN(_31_)
);

NAND2_X1 _82_ (
  .A1(_19_),
  .A2(\fdct_dout[8] ),
  .ZN(_32_)
);

NAND2_X2 _83_ (
  .A1(_31_),
  .A2(_32_),
  .ZN(_07_)
);

NAND2_X4 _84_ (
  .A1(_15_),
  .A2(\dfdct_dout[9] ),
  .ZN(_33_)
);

NAND2_X1 _85_ (
  .A1(_19_),
  .A2(\fdct_dout[9] ),
  .ZN(_34_)
);

NAND2_X2 _86_ (
  .A1(_33_),
  .A2(_34_),
  .ZN(_08_)
);

NAND2_X4 _87_ (
  .A1(_15_),
  .A2(\dfdct_dout[10] ),
  .ZN(_35_)
);

NAND2_X1 _88_ (
  .A1(_19_),
  .A2(\fdct_dout[10] ),
  .ZN(_36_)
);

NAND2_X2 _89_ (
  .A1(_35_),
  .A2(_36_),
  .ZN(_09_)
);

NAND2_X1 _90_ (
  .A1(_14_),
  .A2(\dfdct_dout[11] ),
  .ZN(_37_)
);

NAND2_X1 _91_ (
  .A1(_19_),
  .A2(\fdct_dout[11] ),
  .ZN(_38_)
);

NAND2_X1 _92_ (
  .A1(_37_),
  .A2(_38_),
  .ZN(_10_)
);

NAND2_X1 _93_ (
  .A1(_14_),
  .A2(dc_diff_doe),
  .ZN(_39_)
);

NAND2_X1 _94_ (
  .A1(_19_),
  .A2(qnr_doe),
  .ZN(_40_)
);

NAND2_X1 _95_ (
  .A1(_39_),
  .A2(_40_),
  .ZN(_11_)
);

NAND2_X4 _96_ (
  .A1(_15_),
  .A2(\dfdct_dout[1] ),
  .ZN(_41_)
);

NAND2_X1 _97_ (
  .A1(_13_),
  .A2(\fdct_dout[1] ),
  .ZN(_42_)
);

NAND2_X4 _98_ (
  .A1(_41_),
  .A2(_42_),
  .ZN(_12_)
);

DFF_X1 dc_diff_doe$_DFFE_PP_ (
  .D(_11_),
  .CK(clk),
  .Q(dc_diff_doe),
  .QN(_44_)
);

DFF_X1 \dfdct_dout[0]$_DFFE_PP_  (
  .D(_00_),
  .CK(clk),
  .Q(\dfdct_dout[0] ),
  .QN(_55_)
);

DFF_X1 \dfdct_dout[10]$_DFFE_PP_  (
  .D(_09_),
  .CK(clk),
  .Q(\dfdct_dout[10] ),
  .QN(_46_)
);

DFF_X1 \dfdct_dout[11]$_DFFE_PP_  (
  .D(_10_),
  .CK(clk),
  .Q(\dfdct_dout[11] ),
  .QN(_45_)
);

DFF_X1 \dfdct_dout[1]$_DFFE_PP_  (
  .D(_12_),
  .CK(clk),
  .Q(\dfdct_dout[1] ),
  .QN(_43_)
);

DFF_X1 \dfdct_dout[2]$_DFFE_PP_  (
  .D(_01_),
  .CK(clk),
  .Q(\dfdct_dout[2] ),
  .QN(_54_)
);

DFF_X1 \dfdct_dout[3]$_DFFE_PP_  (
  .D(_02_),
  .CK(clk),
  .Q(\dfdct_dout[3] ),
  .QN(_53_)
);

DFF_X1 \dfdct_dout[4]$_DFFE_PP_  (
  .D(_03_),
  .CK(clk),
  .Q(\dfdct_dout[4] ),
  .QN(_52_)
);

DFF_X1 \dfdct_dout[5]$_DFFE_PP_  (
  .D(_04_),
  .CK(clk),
  .Q(\dfdct_dout[5] ),
  .QN(_51_)
);

DFF_X1 \dfdct_dout[6]$_DFFE_PP_  (
  .D(_05_),
  .CK(clk),
  .Q(\dfdct_dout[6] ),
  .QN(_50_)
);

DFF_X1 \dfdct_dout[7]$_DFFE_PP_  (
  .D(_06_),
  .CK(clk),
  .Q(\dfdct_dout[7] ),
  .QN(_49_)
);

DFF_X1 \dfdct_dout[8]$_DFFE_PP_  (
  .D(_07_),
  .CK(clk),
  .Q(\dfdct_dout[8] ),
  .QN(_48_)
);

DFF_X1 \dfdct_dout[9]$_DFFE_PP_  (
  .D(_08_),
  .CK(clk),
  .Q(\dfdct_dout[9] ),
  .QN(_47_)
);

\$paramod$849c8591669cf197b80ef99050b300773b555aae\fdct  fdct_zigzag (
  .clk(clk),
  .ena(ena),
  .rst(rst),
  .dstrb(dstrb),
  .din(din),
  .dout({\fdct_dout[11] , \fdct_dout[10] , \fdct_dout[9] , \fdct_dout[8] , \fdct_dout[7] , \fdct_dout[6] , \fdct_dout[5] , \fdct_dout[4] , \fdct_dout[3] , \fdct_dout[2] , \fdct_dout[1] , \fdct_dout[0] }),
  .douten(fdct_doe)
);

jpeg_qnr qnr (
  .clk(clk),
  .ena(ena),
  .rst(rst),
  .dstrb(fdct_doe),
  .din({\dfdct_dout[11] , \dfdct_dout[10] , \dfdct_dout[9] , \dfdct_dout[8] , \dfdct_dout[7] , \dfdct_dout[6] , \dfdct_dout[5] , \dfdct_dout[4] , \dfdct_dout[3] , \dfdct_dout[2] , \dfdct_dout[1] , \dfdct_dout[0] }),
  .qnt_val(qnt_val),
  .qnt_cnt(qnt_cnt),
  .dout({\qnr_dout[10] , \qnr_dout[9] , \qnr_dout[8] , \qnr_dout[7] , \qnr_dout[6] , \qnr_dout[5] , \qnr_dout[4] , \qnr_dout[3] , \qnr_dout[2] , \qnr_dout[1] , \qnr_dout[0] }),
  .douten(qnr_doe)
);

jpeg_rle rle (
  .clk(clk),
  .rst(rst),
  .ena(ena),
  .dstrb(dc_diff_doe),
  .din({\qnr_dout[10] , \qnr_dout[10] , \qnr_dout[9] , \qnr_dout[8] , \qnr_dout[7] , \qnr_dout[6] , \qnr_dout[5] , \qnr_dout[4] , \qnr_dout[3] , \qnr_dout[2] , \qnr_dout[1] , \qnr_dout[0] }),
  .size(size),
  .rlen(rlen),
  .amp(amp),
  .douten(douten)
);
endmodule //jpeg_encoder
